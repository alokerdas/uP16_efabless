magic
tech sky130B
magscale 1 2
timestamp 1657859617
<< metal1 >>
rect 71774 702992 71780 703044
rect 71832 703032 71838 703044
rect 72970 703032 72976 703044
rect 71832 703004 72976 703032
rect 71832 702992 71838 703004
rect 72970 702992 72976 703004
rect 73028 702992 73034 703044
rect 201494 702992 201500 703044
rect 201552 703032 201558 703044
rect 202782 703032 202788 703044
rect 201552 703004 202788 703032
rect 201552 702992 201558 703004
rect 202782 702992 202788 703004
rect 202840 702992 202846 703044
rect 170306 700476 170312 700528
rect 170364 700516 170370 700528
rect 192478 700516 192484 700528
rect 170364 700488 192484 700516
rect 170364 700476 170370 700488
rect 192478 700476 192484 700488
rect 192536 700476 192542 700528
rect 255590 700476 255596 700528
rect 255648 700516 255654 700528
rect 283834 700516 283840 700528
rect 255648 700488 283840 700516
rect 255648 700476 255654 700488
rect 283834 700476 283840 700488
rect 283892 700476 283898 700528
rect 331858 700476 331864 700528
rect 331916 700516 331922 700528
rect 397454 700516 397460 700528
rect 331916 700488 397460 700516
rect 331916 700476 331922 700488
rect 397454 700476 397460 700488
rect 397512 700476 397518 700528
rect 154114 700408 154120 700460
rect 154172 700448 154178 700460
rect 242158 700448 242164 700460
rect 154172 700420 242164 700448
rect 154172 700408 154178 700420
rect 242158 700408 242164 700420
rect 242216 700408 242222 700460
rect 265618 700408 265624 700460
rect 265676 700448 265682 700460
rect 348786 700448 348792 700460
rect 265676 700420 348792 700448
rect 265676 700408 265682 700420
rect 348786 700408 348792 700420
rect 348844 700408 348850 700460
rect 89162 700340 89168 700392
rect 89220 700380 89226 700392
rect 257614 700380 257620 700392
rect 89220 700352 257620 700380
rect 89220 700340 89226 700352
rect 257614 700340 257620 700352
rect 257672 700340 257678 700392
rect 324958 700340 324964 700392
rect 325016 700380 325022 700392
rect 332502 700380 332508 700392
rect 325016 700352 332508 700380
rect 325016 700340 325022 700352
rect 332502 700340 332508 700352
rect 332560 700340 332566 700392
rect 347038 700340 347044 700392
rect 347096 700380 347102 700392
rect 462314 700380 462320 700392
rect 347096 700352 462320 700380
rect 347096 700340 347102 700352
rect 462314 700340 462320 700352
rect 462372 700340 462378 700392
rect 24302 700272 24308 700324
rect 24360 700312 24366 700324
rect 192570 700312 192576 700324
rect 24360 700284 192576 700312
rect 24360 700272 24366 700284
rect 192570 700272 192576 700284
rect 192628 700272 192634 700324
rect 258718 700272 258724 700324
rect 258776 700312 258782 700324
rect 413646 700312 413652 700324
rect 258776 700284 413652 700312
rect 258776 700272 258782 700284
rect 413646 700272 413652 700284
rect 413704 700272 413710 700324
rect 218974 699660 218980 699712
rect 219032 699700 219038 699712
rect 220078 699700 220084 699712
rect 219032 699672 220084 699700
rect 219032 699660 219038 699672
rect 220078 699660 220084 699672
rect 220136 699660 220142 699712
rect 266354 697552 266360 697604
rect 266412 697592 266418 697604
rect 267642 697592 267648 697604
rect 266412 697564 267648 697592
rect 266412 697552 266418 697564
rect 267642 697552 267648 697564
rect 267700 697552 267706 697604
rect 264238 696940 264244 696992
rect 264296 696980 264302 696992
rect 580166 696980 580172 696992
rect 264296 696952 580172 696980
rect 264296 696940 264302 696952
rect 580166 696940 580172 696952
rect 580224 696940 580230 696992
rect 3418 683204 3424 683256
rect 3476 683244 3482 683256
rect 257338 683244 257344 683256
rect 3476 683216 257344 683244
rect 3476 683204 3482 683216
rect 257338 683204 257344 683216
rect 257396 683204 257402 683256
rect 253198 683136 253204 683188
rect 253256 683176 253262 683188
rect 580166 683176 580172 683188
rect 253256 683148 580172 683176
rect 253256 683136 253262 683148
rect 580166 683136 580172 683148
rect 580224 683136 580230 683188
rect 3418 670760 3424 670812
rect 3476 670800 3482 670812
rect 258810 670800 258816 670812
rect 3476 670772 258816 670800
rect 3476 670760 3482 670772
rect 258810 670760 258816 670772
rect 258868 670760 258874 670812
rect 251818 670692 251824 670744
rect 251876 670732 251882 670744
rect 580166 670732 580172 670744
rect 251876 670704 580172 670732
rect 251876 670692 251882 670704
rect 580166 670692 580172 670704
rect 580224 670692 580230 670744
rect 3418 656888 3424 656940
rect 3476 656928 3482 656940
rect 192662 656928 192668 656940
rect 3476 656900 192668 656928
rect 3476 656888 3482 656900
rect 192662 656888 192668 656900
rect 192720 656888 192726 656940
rect 261478 643084 261484 643136
rect 261536 643124 261542 643136
rect 580166 643124 580172 643136
rect 261536 643096 580172 643124
rect 261536 643084 261542 643096
rect 580166 643084 580172 643096
rect 580224 643084 580230 643136
rect 3418 632068 3424 632120
rect 3476 632108 3482 632120
rect 259822 632108 259828 632120
rect 3476 632080 259828 632108
rect 3476 632068 3482 632080
rect 259822 632068 259828 632080
rect 259880 632068 259886 632120
rect 249886 630640 249892 630692
rect 249944 630680 249950 630692
rect 580166 630680 580172 630692
rect 249944 630652 580172 630680
rect 249944 630640 249950 630652
rect 580166 630640 580172 630652
rect 580224 630640 580230 630692
rect 2774 619080 2780 619132
rect 2832 619120 2838 619132
rect 4798 619120 4804 619132
rect 2832 619092 4804 619120
rect 2832 619080 2838 619092
rect 4798 619080 4804 619092
rect 4856 619080 4862 619132
rect 251910 616836 251916 616888
rect 251968 616876 251974 616888
rect 580166 616876 580172 616888
rect 251968 616848 580172 616876
rect 251968 616836 251974 616848
rect 580166 616836 580172 616848
rect 580224 616836 580230 616888
rect 3234 605820 3240 605872
rect 3292 605860 3298 605872
rect 259546 605860 259552 605872
rect 3292 605832 259552 605860
rect 3292 605820 3298 605832
rect 259546 605820 259552 605832
rect 259604 605820 259610 605872
rect 261570 590656 261576 590708
rect 261628 590696 261634 590708
rect 579798 590696 579804 590708
rect 261628 590668 579804 590696
rect 261628 590656 261634 590668
rect 579798 590656 579804 590668
rect 579856 590656 579862 590708
rect 136634 590044 136640 590096
rect 136692 590084 136698 590096
rect 256786 590084 256792 590096
rect 136692 590056 256792 590084
rect 136692 590044 136698 590056
rect 256786 590044 256792 590056
rect 256844 590044 256850 590096
rect 104894 589976 104900 590028
rect 104952 590016 104958 590028
rect 257430 590016 257436 590028
rect 104952 589988 257436 590016
rect 104952 589976 104958 589988
rect 257430 589976 257436 589988
rect 257488 589976 257494 590028
rect 252646 589908 252652 589960
rect 252704 589948 252710 589960
rect 429194 589948 429200 589960
rect 252704 589920 429200 589948
rect 252704 589908 252710 589920
rect 429194 589908 429200 589920
rect 429252 589908 429258 589960
rect 2774 566040 2780 566092
rect 2832 566080 2838 566092
rect 4890 566080 4896 566092
rect 2832 566052 4896 566080
rect 2832 566040 2838 566052
rect 4890 566040 4896 566052
rect 4948 566040 4954 566092
rect 2774 553664 2780 553716
rect 2832 553704 2838 553716
rect 4982 553704 4988 553716
rect 2832 553676 4988 553704
rect 2832 553664 2838 553676
rect 4982 553664 4988 553676
rect 5040 553664 5046 553716
rect 279418 536800 279424 536852
rect 279476 536840 279482 536852
rect 376938 536840 376944 536852
rect 279476 536812 376944 536840
rect 279476 536800 279482 536812
rect 376938 536800 376944 536812
rect 376996 536800 377002 536852
rect 278038 535440 278044 535492
rect 278096 535480 278102 535492
rect 377030 535480 377036 535492
rect 278096 535452 377036 535480
rect 278096 535440 278102 535452
rect 377030 535440 377036 535452
rect 377088 535440 377094 535492
rect 278130 534080 278136 534132
rect 278188 534120 278194 534132
rect 376938 534120 376944 534132
rect 278188 534092 376944 534120
rect 278188 534080 278194 534092
rect 376938 534080 376944 534092
rect 376996 534080 377002 534132
rect 275278 532720 275284 532772
rect 275336 532760 275342 532772
rect 377030 532760 377036 532772
rect 275336 532732 377036 532760
rect 275336 532720 275342 532732
rect 377030 532720 377036 532732
rect 377088 532720 377094 532772
rect 278222 531292 278228 531344
rect 278280 531332 278286 531344
rect 376938 531332 376944 531344
rect 278280 531304 376944 531332
rect 278280 531292 278286 531304
rect 376938 531292 376944 531304
rect 376996 531292 377002 531344
rect 273898 529932 273904 529984
rect 273956 529972 273962 529984
rect 376938 529972 376944 529984
rect 273956 529944 376944 529972
rect 273956 529932 273962 529944
rect 376938 529932 376944 529944
rect 376996 529932 377002 529984
rect 273990 528572 273996 528624
rect 274048 528612 274054 528624
rect 376846 528612 376852 528624
rect 274048 528584 376852 528612
rect 274048 528572 274054 528584
rect 376846 528572 376852 528584
rect 376904 528572 376910 528624
rect 471238 510620 471244 510672
rect 471296 510660 471302 510672
rect 579614 510660 579620 510672
rect 471296 510632 579620 510660
rect 471296 510620 471302 510632
rect 579614 510620 579620 510632
rect 579672 510620 579678 510672
rect 295978 509260 295984 509312
rect 296036 509300 296042 509312
rect 376938 509300 376944 509312
rect 296036 509272 376944 509300
rect 296036 509260 296042 509272
rect 376938 509260 376944 509272
rect 376996 509260 377002 509312
rect 296070 507900 296076 507952
rect 296128 507940 296134 507952
rect 376754 507940 376760 507952
rect 296128 507912 376760 507940
rect 296128 507900 296134 507912
rect 376754 507900 376760 507912
rect 376812 507900 376818 507952
rect 271138 507832 271144 507884
rect 271196 507872 271202 507884
rect 377030 507872 377036 507884
rect 271196 507844 377036 507872
rect 271196 507832 271202 507844
rect 377030 507832 377036 507844
rect 377088 507832 377094 507884
rect 3326 501304 3332 501356
rect 3384 501344 3390 501356
rect 7558 501344 7564 501356
rect 3384 501316 7564 501344
rect 3384 501304 3390 501316
rect 7558 501304 7564 501316
rect 7616 501304 7622 501356
rect 123386 498040 123392 498092
rect 123444 498080 123450 498092
rect 124858 498080 124864 498092
rect 123444 498052 124864 498080
rect 123444 498040 123450 498052
rect 124858 498040 124864 498052
rect 124916 498040 124922 498092
rect 287422 497156 287428 497208
rect 287480 497196 287486 497208
rect 397454 497196 397460 497208
rect 287480 497168 397460 497196
rect 287480 497156 287486 497168
rect 397454 497156 397460 497168
rect 397512 497156 397518 497208
rect 288618 497088 288624 497140
rect 288676 497128 288682 497140
rect 398834 497128 398840 497140
rect 288676 497100 398840 497128
rect 288676 497088 288682 497100
rect 398834 497088 398840 497100
rect 398892 497088 398898 497140
rect 119338 497020 119344 497072
rect 119396 497060 119402 497072
rect 279694 497060 279700 497072
rect 119396 497032 279700 497060
rect 119396 497020 119402 497032
rect 279694 497020 279700 497032
rect 279752 497020 279758 497072
rect 288526 497020 288532 497072
rect 288584 497060 288590 497072
rect 398926 497060 398932 497072
rect 288584 497032 398932 497060
rect 288584 497020 288590 497032
rect 398926 497020 398932 497032
rect 398984 497020 398990 497072
rect 126790 496952 126796 497004
rect 126848 496992 126854 497004
rect 282178 496992 282184 497004
rect 126848 496964 282184 496992
rect 126848 496952 126854 496964
rect 282178 496952 282184 496964
rect 282236 496952 282242 497004
rect 292666 496952 292672 497004
rect 292724 496992 292730 497004
rect 403158 496992 403164 497004
rect 292724 496964 403164 496992
rect 292724 496952 292730 496964
rect 403158 496952 403164 496964
rect 403216 496952 403222 497004
rect 125226 496884 125232 496936
rect 125284 496924 125290 496936
rect 285214 496924 285220 496936
rect 125284 496896 285220 496924
rect 125284 496884 125290 496896
rect 285214 496884 285220 496896
rect 285272 496884 285278 496936
rect 285766 496884 285772 496936
rect 285824 496924 285830 496936
rect 404354 496924 404360 496936
rect 285824 496896 404360 496924
rect 285824 496884 285830 496896
rect 404354 496884 404360 496896
rect 404412 496884 404418 496936
rect 115474 496816 115480 496868
rect 115532 496856 115538 496868
rect 116578 496856 116584 496868
rect 115532 496828 116584 496856
rect 115532 496816 115538 496828
rect 116578 496816 116584 496828
rect 116636 496816 116642 496868
rect 287146 496816 287152 496868
rect 287204 496856 287210 496868
rect 409874 496856 409880 496868
rect 287204 496828 409880 496856
rect 287204 496816 287210 496828
rect 409874 496816 409880 496828
rect 409932 496816 409938 496868
rect 249150 484372 249156 484424
rect 249208 484412 249214 484424
rect 580166 484412 580172 484424
rect 249208 484384 580172 484412
rect 249208 484372 249214 484384
rect 580166 484372 580172 484384
rect 580224 484372 580230 484424
rect 3326 474716 3332 474768
rect 3384 474756 3390 474768
rect 261662 474756 261668 474768
rect 3384 474728 261668 474756
rect 3384 474716 3390 474728
rect 261662 474716 261668 474728
rect 261720 474716 261726 474768
rect 247126 470568 247132 470620
rect 247184 470608 247190 470620
rect 579982 470608 579988 470620
rect 247184 470580 579988 470608
rect 247184 470568 247190 470580
rect 579982 470568 579988 470580
rect 580040 470568 580046 470620
rect 3326 462340 3332 462392
rect 3384 462380 3390 462392
rect 175918 462380 175924 462392
rect 3384 462352 175924 462380
rect 3384 462340 3390 462352
rect 175918 462340 175924 462352
rect 175976 462340 175982 462392
rect 247402 456764 247408 456816
rect 247460 456804 247466 456816
rect 580166 456804 580172 456816
rect 247460 456776 580172 456804
rect 247460 456764 247466 456776
rect 580166 456764 580172 456776
rect 580224 456764 580230 456816
rect 3326 448536 3332 448588
rect 3384 448576 3390 448588
rect 262582 448576 262588 448588
rect 3384 448548 262588 448576
rect 3384 448536 3390 448548
rect 262582 448536 262588 448548
rect 262640 448536 262646 448588
rect 245746 430584 245752 430636
rect 245804 430624 245810 430636
rect 579614 430624 579620 430636
rect 245804 430596 579620 430624
rect 245804 430584 245810 430596
rect 579614 430584 579620 430596
rect 579672 430584 579678 430636
rect 97534 426368 97540 426420
rect 97592 426408 97598 426420
rect 295610 426408 295616 426420
rect 97592 426380 295616 426408
rect 97592 426368 97598 426380
rect 295610 426368 295616 426380
rect 295668 426408 295674 426420
rect 296070 426408 296076 426420
rect 295668 426380 296076 426408
rect 295668 426368 295674 426380
rect 296070 426368 296076 426380
rect 296128 426368 296134 426420
rect 3142 422288 3148 422340
rect 3200 422328 3206 422340
rect 261754 422328 261760 422340
rect 3200 422300 261760 422328
rect 3200 422288 3206 422300
rect 261754 422288 261760 422300
rect 261812 422288 261818 422340
rect 247218 418140 247224 418192
rect 247276 418180 247282 418192
rect 579706 418180 579712 418192
rect 247276 418152 579712 418180
rect 247276 418140 247282 418152
rect 579706 418140 579712 418152
rect 579764 418140 579770 418192
rect 155862 414808 155868 414860
rect 155920 414848 155926 414860
rect 284386 414848 284392 414860
rect 155920 414820 284392 414848
rect 155920 414808 155926 414820
rect 284386 414808 284392 414820
rect 284444 414808 284450 414860
rect 151722 414740 151728 414792
rect 151780 414780 151786 414792
rect 283650 414780 283656 414792
rect 151780 414752 283656 414780
rect 151780 414740 151786 414752
rect 283650 414740 283656 414752
rect 283708 414740 283714 414792
rect 146202 414672 146208 414724
rect 146260 414712 146266 414724
rect 281902 414712 281908 414724
rect 146260 414684 281908 414712
rect 146260 414672 146266 414684
rect 281902 414672 281908 414684
rect 281960 414672 281966 414724
rect 291286 414672 291292 414724
rect 291344 414712 291350 414724
rect 401594 414712 401600 414724
rect 291344 414684 401600 414712
rect 291344 414672 291350 414684
rect 401594 414672 401600 414684
rect 401652 414672 401658 414724
rect 3142 409844 3148 409896
rect 3200 409884 3206 409896
rect 234522 409884 234528 409896
rect 3200 409856 234528 409884
rect 3200 409844 3206 409856
rect 234522 409844 234528 409856
rect 234580 409884 234586 409896
rect 263778 409884 263784 409896
rect 234580 409856 263784 409884
rect 234580 409844 234586 409856
rect 263778 409844 263784 409856
rect 263836 409844 263842 409896
rect 248506 406376 248512 406428
rect 248564 406416 248570 406428
rect 580350 406416 580356 406428
rect 248564 406388 580356 406416
rect 248564 406376 248570 406388
rect 580350 406376 580356 406388
rect 580408 406376 580414 406428
rect 246022 404336 246028 404388
rect 246080 404376 246086 404388
rect 579982 404376 579988 404388
rect 246080 404348 579988 404376
rect 246080 404336 246086 404348
rect 579982 404336 579988 404348
rect 580040 404336 580046 404388
rect 124858 401004 124864 401056
rect 124916 401044 124922 401056
rect 283006 401044 283012 401056
rect 124916 401016 283012 401044
rect 124916 401004 124922 401016
rect 283006 401004 283012 401016
rect 283064 401004 283070 401056
rect 121270 400936 121276 400988
rect 121328 400976 121334 400988
rect 281810 400976 281816 400988
rect 121328 400948 281816 400976
rect 121328 400936 121334 400948
rect 281810 400936 281816 400948
rect 281868 400936 281874 400988
rect 122742 400868 122748 400920
rect 122800 400908 122806 400920
rect 283098 400908 283104 400920
rect 122800 400880 283104 400908
rect 122800 400868 122806 400880
rect 283098 400868 283104 400880
rect 283156 400868 283162 400920
rect 254026 399712 254032 399764
rect 254084 399752 254090 399764
rect 266354 399752 266360 399764
rect 254084 399724 266360 399752
rect 254084 399712 254090 399724
rect 266354 399712 266360 399724
rect 266412 399712 266418 399764
rect 161382 399644 161388 399696
rect 161440 399684 161446 399696
rect 285858 399684 285864 399696
rect 161440 399656 285864 399684
rect 161440 399644 161446 399656
rect 285858 399644 285864 399656
rect 285916 399644 285922 399696
rect 140682 399576 140688 399628
rect 140740 399616 140746 399628
rect 280246 399616 280252 399628
rect 140740 399588 280252 399616
rect 140740 399576 140746 399588
rect 280246 399576 280252 399588
rect 280304 399576 280310 399628
rect 118602 399508 118608 399560
rect 118660 399548 118666 399560
rect 278590 399548 278596 399560
rect 118660 399520 278596 399548
rect 118660 399508 118666 399520
rect 278590 399508 278596 399520
rect 278648 399508 278654 399560
rect 121362 399440 121368 399492
rect 121420 399480 121426 399492
rect 280798 399480 280804 399492
rect 121420 399452 280804 399480
rect 121420 399440 121426 399452
rect 280798 399440 280804 399452
rect 280856 399440 280862 399492
rect 136542 398148 136548 398200
rect 136600 398188 136606 398200
rect 280338 398188 280344 398200
rect 136600 398160 280344 398188
rect 136600 398148 136606 398160
rect 280338 398148 280344 398160
rect 280396 398148 280402 398200
rect 97810 398080 97816 398132
rect 97868 398120 97874 398132
rect 277302 398120 277308 398132
rect 97868 398092 277308 398120
rect 97868 398080 97874 398092
rect 277302 398080 277308 398092
rect 277360 398080 277366 398132
rect 3326 397468 3332 397520
rect 3384 397508 3390 397520
rect 263410 397508 263416 397520
rect 3384 397480 263416 397508
rect 3384 397468 3390 397480
rect 263410 397468 263416 397480
rect 263468 397468 263474 397520
rect 97626 397400 97632 397452
rect 97684 397440 97690 397452
rect 295978 397440 295984 397452
rect 97684 397412 295984 397440
rect 97684 397400 97690 397412
rect 295978 397400 295984 397412
rect 296036 397400 296042 397452
rect 99098 397332 99104 397384
rect 99156 397372 99162 397384
rect 275278 397372 275284 397384
rect 99156 397344 275284 397372
rect 99156 397332 99162 397344
rect 275278 397332 275284 397344
rect 275336 397332 275342 397384
rect 131022 396788 131028 396840
rect 131080 396828 131086 396840
rect 279142 396828 279148 396840
rect 131080 396800 279148 396828
rect 131080 396788 131086 396800
rect 279142 396788 279148 396800
rect 279200 396788 279206 396840
rect 99190 396720 99196 396772
rect 99248 396760 99254 396772
rect 275922 396760 275928 396772
rect 99248 396732 275928 396760
rect 99248 396720 99254 396732
rect 275922 396720 275928 396732
rect 275980 396720 275986 396772
rect 294046 396720 294052 396772
rect 294104 396760 294110 396772
rect 405734 396760 405740 396772
rect 294104 396732 405740 396760
rect 294104 396720 294110 396732
rect 405734 396720 405740 396732
rect 405792 396720 405798 396772
rect 275370 396040 275376 396092
rect 275428 396080 275434 396092
rect 275922 396080 275928 396092
rect 275428 396052 275928 396080
rect 275428 396040 275434 396052
rect 275922 396040 275928 396052
rect 275980 396080 275986 396092
rect 278130 396080 278136 396092
rect 275980 396052 278136 396080
rect 275980 396040 275986 396052
rect 278130 396040 278136 396052
rect 278188 396040 278194 396092
rect 98914 395972 98920 396024
rect 98972 396012 98978 396024
rect 273990 396012 273996 396024
rect 98972 395984 273996 396012
rect 98972 395972 98978 395984
rect 273990 395972 273996 395984
rect 274048 395972 274054 396024
rect 99006 395904 99012 395956
rect 99064 395944 99070 395956
rect 273898 395944 273904 395956
rect 99064 395916 273904 395944
rect 99064 395904 99070 395916
rect 273898 395904 273904 395916
rect 273956 395944 273962 395956
rect 274174 395944 274180 395956
rect 273956 395916 274180 395944
rect 273956 395904 273962 395916
rect 274174 395904 274180 395916
rect 274232 395904 274238 395956
rect 277302 395904 277308 395956
rect 277360 395944 277366 395956
rect 279418 395944 279424 395956
rect 277360 395916 279424 395944
rect 277360 395904 277366 395916
rect 279418 395904 279424 395916
rect 279476 395904 279482 395956
rect 294138 395428 294144 395480
rect 294196 395468 294202 395480
rect 404446 395468 404452 395480
rect 294196 395440 404452 395468
rect 294196 395428 294202 395440
rect 404446 395428 404452 395440
rect 404504 395428 404510 395480
rect 116578 395360 116584 395412
rect 116636 395400 116642 395412
rect 271966 395400 271972 395412
rect 116636 395372 271972 395400
rect 116636 395360 116642 395372
rect 271966 395360 271972 395372
rect 272024 395360 272030 395412
rect 290734 395360 290740 395412
rect 290792 395400 290798 395412
rect 400214 395400 400220 395412
rect 290792 395372 400220 395400
rect 290792 395360 290798 395372
rect 400214 395360 400220 395372
rect 400272 395360 400278 395412
rect 114462 395292 114468 395344
rect 114520 395332 114526 395344
rect 272518 395332 272524 395344
rect 114520 395304 272524 395332
rect 114520 395292 114526 395304
rect 272518 395292 272524 395304
rect 272576 395292 272582 395344
rect 294598 395292 294604 395344
rect 294656 395332 294662 395344
rect 440234 395332 440240 395344
rect 294656 395304 440240 395332
rect 294656 395292 294662 395304
rect 440234 395292 440240 395304
rect 440292 395292 440298 395344
rect 254578 394136 254584 394188
rect 254636 394176 254642 394188
rect 265618 394176 265624 394188
rect 254636 394148 265624 394176
rect 254636 394136 254642 394148
rect 265618 394136 265624 394148
rect 265676 394136 265682 394188
rect 242158 394068 242164 394120
rect 242216 394108 242222 394120
rect 257154 394108 257160 394120
rect 242216 394080 257160 394108
rect 242216 394068 242222 394080
rect 257154 394068 257160 394080
rect 257212 394068 257218 394120
rect 291378 394068 291384 394120
rect 291436 394108 291442 394120
rect 425054 394108 425060 394120
rect 291436 394080 425060 394108
rect 291436 394068 291442 394080
rect 425054 394068 425060 394080
rect 425112 394068 425118 394120
rect 113082 394000 113088 394052
rect 113140 394040 113146 394052
rect 272610 394040 272616 394052
rect 113140 394012 272616 394040
rect 113140 394000 113146 394012
rect 272610 394000 272616 394012
rect 272668 394000 272674 394052
rect 292390 394000 292396 394052
rect 292448 394040 292454 394052
rect 429194 394040 429200 394052
rect 292448 394012 429200 394040
rect 292448 394000 292454 394012
rect 429194 394000 429200 394012
rect 429252 394000 429258 394052
rect 3602 393932 3608 393984
rect 3660 393972 3666 393984
rect 262122 393972 262128 393984
rect 3660 393944 262128 393972
rect 3660 393932 3666 393944
rect 262122 393932 262128 393944
rect 262180 393932 262186 393984
rect 293494 393932 293500 393984
rect 293552 393972 293558 393984
rect 434714 393972 434720 393984
rect 293552 393944 434720 393972
rect 293552 393932 293558 393944
rect 434714 393932 434720 393944
rect 434772 393932 434778 393984
rect 260466 393428 260472 393440
rect 238726 393400 260472 393428
rect 233786 393320 233792 393372
rect 233844 393360 233850 393372
rect 238726 393360 238754 393400
rect 260466 393388 260472 393400
rect 260524 393388 260530 393440
rect 233844 393332 238754 393360
rect 233844 393320 233850 393332
rect 252922 393320 252928 393372
rect 252980 393360 252986 393372
rect 258718 393360 258724 393372
rect 252980 393332 258724 393360
rect 252980 393320 252986 393332
rect 258718 393320 258724 393332
rect 258776 393320 258782 393372
rect 220078 392844 220084 392896
rect 220136 392884 220142 392896
rect 256234 392884 256240 392896
rect 220136 392856 256240 392884
rect 220136 392844 220142 392856
rect 256234 392844 256240 392856
rect 256292 392844 256298 392896
rect 253014 392776 253020 392828
rect 253072 392816 253078 392828
rect 477494 392816 477500 392828
rect 253072 392788 477500 392816
rect 253072 392776 253078 392788
rect 477494 392776 477500 392788
rect 477552 392776 477558 392828
rect 7558 392708 7564 392760
rect 7616 392748 7622 392760
rect 261938 392748 261944 392760
rect 7616 392720 261944 392748
rect 7616 392708 7622 392720
rect 261938 392708 261944 392720
rect 261996 392708 262002 392760
rect 251266 392640 251272 392692
rect 251324 392680 251330 392692
rect 542354 392680 542360 392692
rect 251324 392652 542360 392680
rect 251324 392640 251330 392652
rect 542354 392640 542360 392652
rect 542412 392640 542418 392692
rect 192570 392572 192576 392624
rect 192628 392612 192634 392624
rect 233970 392612 233976 392624
rect 192628 392584 233976 392612
rect 192628 392572 192634 392584
rect 233970 392572 233976 392584
rect 234028 392572 234034 392624
rect 248782 392572 248788 392624
rect 248840 392612 248846 392624
rect 580534 392612 580540 392624
rect 248840 392584 580540 392612
rect 248840 392572 248846 392584
rect 580534 392572 580540 392584
rect 580592 392572 580598 392624
rect 248506 392436 248512 392488
rect 248564 392476 248570 392488
rect 249610 392476 249616 392488
rect 248564 392448 249616 392476
rect 248564 392436 248570 392448
rect 249610 392436 249616 392448
rect 249668 392436 249674 392488
rect 233970 391960 233976 392012
rect 234028 392000 234034 392012
rect 258718 392000 258724 392012
rect 234028 391972 258724 392000
rect 234028 391960 234034 391972
rect 258718 391960 258724 391972
rect 258776 391960 258782 392012
rect 192662 391552 192668 391604
rect 192720 391592 192726 391604
rect 259270 391592 259276 391604
rect 192720 391564 259276 391592
rect 192720 391552 192726 391564
rect 259270 391552 259276 391564
rect 259328 391552 259334 391604
rect 254394 391484 254400 391536
rect 254452 391524 254458 391536
rect 324958 391524 324964 391536
rect 254452 391496 324964 391524
rect 254452 391484 254458 391496
rect 324958 391484 324964 391496
rect 325016 391484 325022 391536
rect 253474 391416 253480 391468
rect 253532 391456 253538 391468
rect 331858 391456 331864 391468
rect 253532 391428 331864 391456
rect 253532 391416 253538 391428
rect 331858 391416 331864 391428
rect 331916 391416 331922 391468
rect 252738 391348 252744 391400
rect 252796 391388 252802 391400
rect 347038 391388 347044 391400
rect 252796 391360 347044 391388
rect 252796 391348 252802 391360
rect 347038 391348 347044 391360
rect 347096 391348 347102 391400
rect 6914 391280 6920 391332
rect 6972 391320 6978 391332
rect 258534 391320 258540 391332
rect 6972 391292 258540 391320
rect 6972 391280 6978 391292
rect 258534 391280 258540 391292
rect 258592 391280 258598 391332
rect 4982 391212 4988 391264
rect 5040 391252 5046 391264
rect 260926 391252 260932 391264
rect 5040 391224 260932 391252
rect 5040 391212 5046 391224
rect 260926 391212 260932 391224
rect 260984 391212 260990 391264
rect 251358 390532 251364 390584
rect 251416 390572 251422 390584
rect 253198 390572 253204 390584
rect 251416 390544 253204 390572
rect 251416 390532 251422 390544
rect 253198 390532 253204 390544
rect 253256 390532 253262 390584
rect 258810 390532 258816 390584
rect 258868 390572 258874 390584
rect 260190 390572 260196 390584
rect 258868 390544 260196 390572
rect 258868 390532 258874 390544
rect 260190 390532 260196 390544
rect 260248 390532 260254 390584
rect 273070 390464 273076 390516
rect 273128 390504 273134 390516
rect 394694 390504 394700 390516
rect 273128 390476 394700 390504
rect 273128 390464 273134 390476
rect 394694 390464 394700 390476
rect 394752 390464 394758 390516
rect 250162 390124 250168 390176
rect 250220 390164 250226 390176
rect 261478 390164 261484 390176
rect 250220 390136 261484 390164
rect 250220 390124 250226 390136
rect 261478 390124 261484 390136
rect 261536 390124 261542 390176
rect 249334 390056 249340 390108
rect 249392 390096 249398 390108
rect 261570 390096 261576 390108
rect 249392 390068 261576 390096
rect 249392 390056 249398 390068
rect 261570 390056 261576 390068
rect 261628 390056 261634 390108
rect 250990 389988 250996 390040
rect 251048 390028 251054 390040
rect 264238 390028 264244 390040
rect 251048 390000 264244 390028
rect 251048 389988 251054 390000
rect 264238 389988 264244 390000
rect 264296 389988 264302 390040
rect 271966 389988 271972 390040
rect 272024 390028 272030 390040
rect 273070 390028 273076 390040
rect 272024 390000 273076 390028
rect 272024 389988 272030 390000
rect 273070 389988 273076 390000
rect 273128 389988 273134 390040
rect 71774 389920 71780 389972
rect 71832 389960 71838 389972
rect 257614 389960 257620 389972
rect 71832 389932 257620 389960
rect 71832 389920 71838 389932
rect 257614 389920 257620 389932
rect 257672 389920 257678 389972
rect 252002 389852 252008 389904
rect 252060 389892 252066 389904
rect 527174 389892 527180 389904
rect 252060 389864 527180 389892
rect 252060 389852 252066 389864
rect 527174 389852 527180 389864
rect 527232 389852 527238 389904
rect 248414 389784 248420 389836
rect 248472 389824 248478 389836
rect 580442 389824 580448 389836
rect 248472 389796 580448 389824
rect 248472 389784 248478 389796
rect 580442 389784 580448 389796
rect 580500 389784 580506 389836
rect 287146 389716 287152 389768
rect 287204 389756 287210 389768
rect 287974 389756 287980 389768
rect 287204 389728 287980 389756
rect 287204 389716 287210 389728
rect 287974 389716 287980 389728
rect 288032 389716 288038 389768
rect 288526 389308 288532 389360
rect 288584 389348 288590 389360
rect 289630 389348 289636 389360
rect 288584 389320 289636 389348
rect 288584 389308 288590 389320
rect 289630 389308 289636 389320
rect 289688 389308 289694 389360
rect 254946 388832 254952 388884
rect 255004 388872 255010 388884
rect 299474 388872 299480 388884
rect 255004 388844 299480 388872
rect 255004 388832 255010 388844
rect 299474 388832 299480 388844
rect 299532 388832 299538 388884
rect 201494 388764 201500 388816
rect 201552 388804 201558 388816
rect 255958 388804 255964 388816
rect 201552 388776 255964 388804
rect 201552 388764 201558 388776
rect 255958 388764 255964 388776
rect 256016 388764 256022 388816
rect 254302 388696 254308 388748
rect 254360 388736 254366 388748
rect 364334 388736 364340 388748
rect 254360 388708 364340 388736
rect 254360 388696 254366 388708
rect 364334 388696 364340 388708
rect 364392 388696 364398 388748
rect 40034 388628 40040 388680
rect 40092 388668 40098 388680
rect 258166 388668 258172 388680
rect 40092 388640 258172 388668
rect 40092 388628 40098 388640
rect 258166 388628 258172 388640
rect 258224 388628 258230 388680
rect 252462 388560 252468 388612
rect 252520 388600 252526 388612
rect 494054 388600 494060 388612
rect 252520 388572 494060 388600
rect 252520 388560 252526 388572
rect 494054 388560 494060 388572
rect 494112 388560 494118 388612
rect 4890 388492 4896 388544
rect 4948 388532 4954 388544
rect 261294 388532 261300 388544
rect 4948 388504 261300 388532
rect 4948 388492 4954 388504
rect 261294 388492 261300 388504
rect 261352 388492 261358 388544
rect 3510 388424 3516 388476
rect 3568 388464 3574 388476
rect 261478 388464 261484 388476
rect 3568 388436 261484 388464
rect 3568 388424 3574 388436
rect 261478 388424 261484 388436
rect 261536 388424 261542 388476
rect 283006 388424 283012 388476
rect 283064 388464 283070 388476
rect 284110 388464 284116 388476
rect 283064 388436 284116 388464
rect 283064 388424 283070 388436
rect 284110 388424 284116 388436
rect 284168 388424 284174 388476
rect 285766 388424 285772 388476
rect 285824 388464 285830 388476
rect 286870 388464 286876 388476
rect 285824 388436 286876 388464
rect 285824 388424 285830 388436
rect 286870 388424 286876 388436
rect 286928 388424 286934 388476
rect 294046 388424 294052 388476
rect 294104 388464 294110 388476
rect 295150 388464 295156 388476
rect 294104 388436 295156 388464
rect 294104 388424 294110 388436
rect 295150 388424 295156 388436
rect 295208 388424 295214 388476
rect 419534 388464 419540 388476
rect 296686 388436 419540 388464
rect 290182 388356 290188 388408
rect 290240 388396 290246 388408
rect 296686 388396 296714 388436
rect 419534 388424 419540 388436
rect 419592 388424 419598 388476
rect 290240 388368 296714 388396
rect 290240 388356 290246 388368
rect 234614 387404 234620 387456
rect 234672 387444 234678 387456
rect 255682 387444 255688 387456
rect 234672 387416 255688 387444
rect 234672 387404 234678 387416
rect 255682 387404 255688 387416
rect 255740 387404 255746 387456
rect 192478 387336 192484 387388
rect 192536 387376 192542 387388
rect 256510 387376 256516 387388
rect 192536 387348 256516 387376
rect 192536 387336 192542 387348
rect 256510 387336 256516 387348
rect 256568 387336 256574 387388
rect 248322 387268 248328 387320
rect 248380 387308 248386 387320
rect 471238 387308 471244 387320
rect 248380 387280 471244 387308
rect 248380 387268 248386 387280
rect 471238 387268 471244 387280
rect 471296 387268 471302 387320
rect 3418 387200 3424 387252
rect 3476 387240 3482 387252
rect 260650 387240 260656 387252
rect 3476 387212 260656 387240
rect 3476 387200 3482 387212
rect 260650 387200 260656 387212
rect 260708 387200 260714 387252
rect 251634 387132 251640 387184
rect 251692 387172 251698 387184
rect 558914 387172 558920 387184
rect 251692 387144 558920 387172
rect 251692 387132 251698 387144
rect 558914 387132 558920 387144
rect 558972 387132 558978 387184
rect 249242 387064 249248 387116
rect 249300 387104 249306 387116
rect 580258 387104 580264 387116
rect 249300 387076 580264 387104
rect 249300 387064 249306 387076
rect 580258 387064 580264 387076
rect 580316 387064 580322 387116
rect 249978 386520 249984 386572
rect 250036 386560 250042 386572
rect 251910 386560 251916 386572
rect 250036 386532 251916 386560
rect 250036 386520 250042 386532
rect 251910 386520 251916 386532
rect 251968 386520 251974 386572
rect 261754 386520 261760 386572
rect 261812 386560 261818 386572
rect 263134 386560 263140 386572
rect 261812 386532 263140 386560
rect 261812 386520 261818 386532
rect 263134 386520 263140 386532
rect 263192 386520 263198 386572
rect 247770 386452 247776 386504
rect 247828 386492 247834 386504
rect 249150 386492 249156 386504
rect 247828 386464 249156 386492
rect 247828 386452 247834 386464
rect 249150 386452 249156 386464
rect 249208 386452 249214 386504
rect 250806 386452 250812 386504
rect 250864 386492 250870 386504
rect 251818 386492 251824 386504
rect 250864 386464 251824 386492
rect 250864 386452 250870 386464
rect 251818 386452 251824 386464
rect 251876 386452 251882 386504
rect 257338 386452 257344 386504
rect 257396 386492 257402 386504
rect 258994 386492 259000 386504
rect 257396 386464 259000 386492
rect 257396 386452 257402 386464
rect 258994 386452 259000 386464
rect 259052 386452 259058 386504
rect 261662 386452 261668 386504
rect 261720 386492 261726 386504
rect 262306 386492 262312 386504
rect 261720 386464 262312 386492
rect 261720 386452 261726 386464
rect 262306 386452 262312 386464
rect 262364 386452 262370 386504
rect 281626 386492 281632 386504
rect 273226 386464 281632 386492
rect 235810 386384 235816 386436
rect 235868 386424 235874 386436
rect 273226 386424 273254 386464
rect 281626 386452 281632 386464
rect 281684 386452 281690 386504
rect 235868 386396 273254 386424
rect 235868 386384 235874 386396
rect 275370 386384 275376 386436
rect 275428 386424 275434 386436
rect 275830 386424 275836 386436
rect 275428 386396 275836 386424
rect 275428 386384 275434 386396
rect 275830 386384 275836 386396
rect 275888 386384 275894 386436
rect 97718 386316 97724 386368
rect 97776 386356 97782 386368
rect 271506 386356 271512 386368
rect 97776 386328 271512 386356
rect 97776 386316 97782 386328
rect 271506 386316 271512 386328
rect 271564 386316 271570 386368
rect 393314 386356 393320 386368
rect 273226 386328 393320 386356
rect 272518 386248 272524 386300
rect 272576 386288 272582 386300
rect 272794 386288 272800 386300
rect 272576 386260 272800 386288
rect 272576 386248 272582 386260
rect 272794 386248 272800 386260
rect 272852 386288 272858 386300
rect 273226 386288 273254 386328
rect 393314 386316 393320 386328
rect 393372 386316 393378 386368
rect 391934 386288 391940 386300
rect 272852 386260 273254 386288
rect 287026 386260 391940 386288
rect 272852 386248 272858 386260
rect 272242 386180 272248 386232
rect 272300 386220 272306 386232
rect 272610 386220 272616 386232
rect 272300 386192 272616 386220
rect 272300 386180 272306 386192
rect 272610 386180 272616 386192
rect 272668 386220 272674 386232
rect 287026 386220 287054 386260
rect 391934 386248 391940 386260
rect 391992 386248 391998 386300
rect 272668 386192 287054 386220
rect 272668 386180 272674 386192
rect 175918 385840 175924 385892
rect 175976 385880 175982 385892
rect 235534 385880 235540 385892
rect 175976 385852 235540 385880
rect 175976 385840 175982 385852
rect 235534 385840 235540 385852
rect 235592 385840 235598 385892
rect 125502 385772 125508 385824
rect 125560 385812 125566 385824
rect 278130 385812 278136 385824
rect 125560 385784 278136 385812
rect 125560 385772 125566 385784
rect 278130 385772 278136 385784
rect 278188 385772 278194 385824
rect 99282 385704 99288 385756
rect 99340 385744 99346 385756
rect 274818 385744 274824 385756
rect 99340 385716 274824 385744
rect 99340 385704 99346 385716
rect 274818 385704 274824 385716
rect 274876 385744 274882 385756
rect 278222 385744 278228 385756
rect 274876 385716 278228 385744
rect 274876 385704 274882 385716
rect 278222 385704 278228 385716
rect 278280 385704 278286 385756
rect 97902 385636 97908 385688
rect 97960 385676 97966 385688
rect 276474 385676 276480 385688
rect 97960 385648 276480 385676
rect 97960 385636 97966 385648
rect 276474 385636 276480 385648
rect 276532 385676 276538 385688
rect 278038 385676 278044 385688
rect 276532 385648 278044 385676
rect 276532 385636 276538 385648
rect 278038 385636 278044 385648
rect 278096 385636 278102 385688
rect 289262 385636 289268 385688
rect 289320 385676 289326 385688
rect 415394 385676 415400 385688
rect 289320 385648 415400 385676
rect 289320 385636 289326 385648
rect 415394 385636 415400 385648
rect 415452 385636 415458 385688
rect 244918 385296 244924 385348
rect 244976 385336 244982 385348
rect 253842 385336 253848 385348
rect 244976 385308 253848 385336
rect 244976 385296 244982 385308
rect 253842 385296 253848 385308
rect 253900 385296 253906 385348
rect 247126 385228 247132 385280
rect 247184 385268 247190 385280
rect 247954 385268 247960 385280
rect 247184 385240 247960 385268
rect 247184 385228 247190 385240
rect 247954 385228 247960 385240
rect 248012 385228 248018 385280
rect 251266 385228 251272 385280
rect 251324 385268 251330 385280
rect 252094 385268 252100 385280
rect 251324 385240 252100 385268
rect 251324 385228 251330 385240
rect 252094 385228 252100 385240
rect 252152 385228 252158 385280
rect 252646 385228 252652 385280
rect 252704 385268 252710 385280
rect 253198 385268 253204 385280
rect 252704 385240 253204 385268
rect 252704 385228 252710 385240
rect 253198 385228 253204 385240
rect 253256 385228 253262 385280
rect 262858 385268 262864 385280
rect 253906 385240 262864 385268
rect 235534 385160 235540 385212
rect 235592 385200 235598 385212
rect 235718 385200 235724 385212
rect 235592 385172 235724 385200
rect 235592 385160 235598 385172
rect 235718 385160 235724 385172
rect 235776 385200 235782 385212
rect 253906 385200 253934 385240
rect 262858 385228 262864 385240
rect 262916 385228 262922 385280
rect 235776 385172 253934 385200
rect 235776 385160 235782 385172
rect 254026 385160 254032 385212
rect 254084 385200 254090 385212
rect 255130 385200 255136 385212
rect 254084 385172 255136 385200
rect 254084 385160 254090 385172
rect 255130 385160 255136 385172
rect 255188 385160 255194 385212
rect 259546 385160 259552 385212
rect 259604 385200 259610 385212
rect 260098 385200 260104 385212
rect 259604 385172 260104 385200
rect 259604 385160 259610 385172
rect 260098 385160 260104 385172
rect 260156 385160 260162 385212
rect 280246 385160 280252 385212
rect 280304 385200 280310 385212
rect 281350 385200 281356 385212
rect 280304 385172 281356 385200
rect 280304 385160 280310 385172
rect 281350 385160 281356 385172
rect 281408 385160 281414 385212
rect 252922 385092 252928 385144
rect 252980 385132 252986 385144
rect 253750 385132 253756 385144
rect 252980 385104 253756 385132
rect 252980 385092 252986 385104
rect 253750 385092 253756 385104
rect 253808 385092 253814 385144
rect 253842 385092 253848 385144
rect 253900 385132 253906 385144
rect 577958 385132 577964 385144
rect 253900 385104 577964 385132
rect 253900 385092 253906 385104
rect 577958 385092 577964 385104
rect 578016 385092 578022 385144
rect 244090 385024 244096 385076
rect 244148 385064 244154 385076
rect 577774 385064 577780 385076
rect 244148 385036 577780 385064
rect 244148 385024 244154 385036
rect 577774 385024 577780 385036
rect 577832 385024 577838 385076
rect 282178 384956 282184 385008
rect 282236 384996 282242 385008
rect 286318 384996 286324 385008
rect 282236 384968 286324 384996
rect 282236 384956 282242 384968
rect 286318 384956 286324 384968
rect 286376 384956 286382 385008
rect 241054 384820 241060 384872
rect 241112 384860 241118 384872
rect 295334 384860 295340 384872
rect 241112 384832 295340 384860
rect 241112 384820 241118 384832
rect 295334 384820 295340 384832
rect 295392 384820 295398 384872
rect 236822 384752 236828 384804
rect 236880 384792 236886 384804
rect 266998 384792 267004 384804
rect 236880 384764 267004 384792
rect 236880 384752 236886 384764
rect 266998 384752 267004 384764
rect 267056 384752 267062 384804
rect 286778 384752 286784 384804
rect 286836 384792 286842 384804
rect 296806 384792 296812 384804
rect 286836 384764 296812 384792
rect 286836 384752 286842 384764
rect 296806 384752 296812 384764
rect 296864 384752 296870 384804
rect 246390 384684 246396 384736
rect 246448 384724 246454 384736
rect 293770 384724 293776 384736
rect 246448 384696 293776 384724
rect 246448 384684 246454 384696
rect 293770 384684 293776 384696
rect 293828 384684 293834 384736
rect 174538 384616 174544 384668
rect 174596 384656 174602 384668
rect 270310 384656 270316 384668
rect 174596 384628 270316 384656
rect 174596 384616 174602 384628
rect 270310 384616 270316 384628
rect 270368 384616 270374 384668
rect 285582 384616 285588 384668
rect 285640 384656 285646 384668
rect 301866 384656 301872 384668
rect 285640 384628 301872 384656
rect 285640 384616 285646 384628
rect 301866 384616 301872 384628
rect 301924 384616 301930 384668
rect 243814 384548 243820 384600
rect 243872 384588 243878 384600
rect 579982 384588 579988 384600
rect 243872 384560 579988 384588
rect 243872 384548 243878 384560
rect 579982 384548 579988 384560
rect 580040 384548 580046 384600
rect 242802 384480 242808 384532
rect 242860 384520 242866 384532
rect 580534 384520 580540 384532
rect 242860 384492 580540 384520
rect 242860 384480 242866 384492
rect 580534 384480 580540 384492
rect 580592 384480 580598 384532
rect 267642 384412 267648 384464
rect 267700 384452 267706 384464
rect 291838 384452 291844 384464
rect 267700 384424 291844 384452
rect 267700 384412 267706 384424
rect 291838 384412 291844 384424
rect 291896 384412 291902 384464
rect 235626 384344 235632 384396
rect 235684 384384 235690 384396
rect 269758 384384 269764 384396
rect 235684 384356 269764 384384
rect 235684 384344 235690 384356
rect 269758 384344 269764 384356
rect 269816 384344 269822 384396
rect 264882 384276 264888 384328
rect 264940 384316 264946 384328
rect 301774 384316 301780 384328
rect 264940 384288 301780 384316
rect 264940 384276 264946 384288
rect 301774 384276 301780 384288
rect 301832 384276 301838 384328
rect 231118 384208 231124 384260
rect 231176 384248 231182 384260
rect 269482 384248 269488 384260
rect 231176 384220 269488 384248
rect 231176 384208 231182 384220
rect 269482 384208 269488 384220
rect 269540 384208 269546 384260
rect 279510 384208 279516 384260
rect 279568 384248 279574 384260
rect 344646 384248 344652 384260
rect 279568 384220 344652 384248
rect 279568 384208 279574 384220
rect 344646 384208 344652 384220
rect 344704 384208 344710 384260
rect 274450 384140 274456 384192
rect 274508 384180 274514 384192
rect 300118 384180 300124 384192
rect 274508 384152 300124 384180
rect 274508 384140 274514 384152
rect 300118 384140 300124 384152
rect 300176 384140 300182 384192
rect 241330 384072 241336 384124
rect 241388 384112 241394 384124
rect 289722 384112 289728 384124
rect 241388 384084 289728 384112
rect 241388 384072 241394 384084
rect 289722 384072 289728 384084
rect 289780 384072 289786 384124
rect 291286 384072 291292 384124
rect 291344 384112 291350 384124
rect 291838 384112 291844 384124
rect 291344 384084 291844 384112
rect 291344 384072 291350 384084
rect 291838 384072 291844 384084
rect 291896 384072 291902 384124
rect 300486 384112 300492 384124
rect 291948 384084 300492 384112
rect 240042 384004 240048 384056
rect 240100 384044 240106 384056
rect 290918 384044 290924 384056
rect 240100 384016 290924 384044
rect 240100 384004 240106 384016
rect 290918 384004 290924 384016
rect 290976 384004 290982 384056
rect 291746 384004 291752 384056
rect 291804 384044 291810 384056
rect 291948 384044 291976 384084
rect 300486 384072 300492 384084
rect 300544 384072 300550 384124
rect 291804 384016 291976 384044
rect 291804 384004 291810 384016
rect 296530 384004 296536 384056
rect 296588 384044 296594 384056
rect 344278 384044 344284 384056
rect 296588 384016 344284 384044
rect 296588 384004 296594 384016
rect 344278 384004 344284 384016
rect 344336 384004 344342 384056
rect 233970 383936 233976 383988
rect 234028 383976 234034 383988
rect 275554 383976 275560 383988
rect 234028 383948 275560 383976
rect 234028 383936 234034 383948
rect 275554 383936 275560 383948
rect 275612 383936 275618 383988
rect 293402 383936 293408 383988
rect 293460 383976 293466 383988
rect 344094 383976 344100 383988
rect 293460 383948 344100 383976
rect 293460 383936 293466 383948
rect 344094 383936 344100 383948
rect 344152 383936 344158 383988
rect 248874 383868 248880 383920
rect 248932 383908 248938 383920
rect 264514 383908 264520 383920
rect 248932 383880 264520 383908
rect 248932 383868 248938 383880
rect 264514 383868 264520 383880
rect 264572 383868 264578 383920
rect 285122 383868 285128 383920
rect 285180 383908 285186 383920
rect 347774 383908 347780 383920
rect 285180 383880 347780 383908
rect 285180 383868 285186 383880
rect 347774 383868 347780 383880
rect 347832 383868 347838 383920
rect 245194 383800 245200 383852
rect 245252 383840 245258 383852
rect 261202 383840 261208 383852
rect 245252 383812 261208 383840
rect 245252 383800 245258 383812
rect 261202 383800 261208 383812
rect 261260 383800 261266 383852
rect 290642 383800 290648 383852
rect 290700 383840 290706 383852
rect 300210 383840 300216 383852
rect 290700 383812 300216 383840
rect 290700 383800 290706 383812
rect 300210 383800 300216 383812
rect 300268 383800 300274 383852
rect 239398 383732 239404 383784
rect 239456 383772 239462 383784
rect 270034 383772 270040 383784
rect 239456 383744 270040 383772
rect 239456 383732 239462 383744
rect 270034 383732 270040 383744
rect 270092 383732 270098 383784
rect 292758 383732 292764 383784
rect 292816 383772 292822 383784
rect 301498 383772 301504 383784
rect 292816 383744 301504 383772
rect 292816 383732 292822 383744
rect 301498 383732 301504 383744
rect 301556 383732 301562 383784
rect 261294 383664 261300 383716
rect 261352 383704 261358 383716
rect 274542 383704 274548 383716
rect 261352 383676 274548 383704
rect 261352 383664 261358 383676
rect 274542 383664 274548 383676
rect 274600 383664 274606 383716
rect 283558 383664 283564 383716
rect 283616 383704 283622 383716
rect 291102 383704 291108 383716
rect 283616 383676 291108 383704
rect 283616 383664 283622 383676
rect 291102 383664 291108 383676
rect 291160 383664 291166 383716
rect 294506 383664 294512 383716
rect 294564 383704 294570 383716
rect 300394 383704 300400 383716
rect 294564 383676 300400 383704
rect 294564 383664 294570 383676
rect 300394 383664 300400 383676
rect 300452 383664 300458 383716
rect 245654 383256 245660 383308
rect 245712 383296 245718 383308
rect 248874 383296 248880 383308
rect 245712 383268 248880 383296
rect 245712 383256 245718 383268
rect 248874 383256 248880 383268
rect 248932 383256 248938 383308
rect 244642 383188 244648 383240
rect 244700 383228 244706 383240
rect 244700 383200 248644 383228
rect 244700 383188 244706 383200
rect 245470 383120 245476 383172
rect 245528 383160 245534 383172
rect 248616 383160 248644 383200
rect 249058 383188 249064 383240
rect 249116 383228 249122 383240
rect 577590 383228 577596 383240
rect 249116 383200 577596 383228
rect 249116 383188 249122 383200
rect 577590 383188 577596 383200
rect 577648 383188 577654 383240
rect 578050 383160 578056 383172
rect 245528 383132 248552 383160
rect 248616 383132 578056 383160
rect 245528 383120 245534 383132
rect 235442 383052 235448 383104
rect 235500 383092 235506 383104
rect 248524 383092 248552 383132
rect 578050 383120 578056 383132
rect 578108 383120 578114 383172
rect 580258 383092 580264 383104
rect 235500 383064 245792 383092
rect 248524 383064 580264 383092
rect 235500 383052 235506 383064
rect 245764 383024 245792 383064
rect 580258 383052 580264 383064
rect 580316 383052 580322 383104
rect 264790 383024 264796 383036
rect 245764 382996 264796 383024
rect 264790 382984 264796 382996
rect 264848 382984 264854 383036
rect 3786 382916 3792 382968
rect 3844 382956 3850 382968
rect 245654 382956 245660 382968
rect 3844 382928 245660 382956
rect 3844 382916 3850 382928
rect 245654 382916 245660 382928
rect 245712 382916 245718 382968
rect 245746 382916 245752 382968
rect 245804 382956 245810 382968
rect 246850 382956 246856 382968
rect 245804 382928 246856 382956
rect 245804 382916 245810 382928
rect 246850 382916 246856 382928
rect 246908 382916 246914 382968
rect 258626 382916 258632 382968
rect 258684 382956 258690 382968
rect 264054 382956 264060 382968
rect 258684 382928 264060 382956
rect 258684 382916 258690 382928
rect 264054 382916 264060 382928
rect 264112 382956 264118 382968
rect 264882 382956 264888 382968
rect 264112 382928 264888 382956
rect 264112 382916 264118 382928
rect 264882 382916 264888 382928
rect 264940 382916 264946 382968
rect 291102 382916 291108 382968
rect 291160 382956 291166 382968
rect 322934 382956 322940 382968
rect 291160 382928 322940 382956
rect 291160 382916 291166 382928
rect 322934 382916 322940 382928
rect 322992 382916 322998 382968
rect 235166 382848 235172 382900
rect 235224 382888 235230 382900
rect 264238 382888 264244 382900
rect 235224 382860 264244 382888
rect 235224 382848 235230 382860
rect 264238 382848 264244 382860
rect 264296 382848 264302 382900
rect 234154 382780 234160 382832
rect 234212 382820 234218 382832
rect 275002 382820 275008 382832
rect 234212 382792 275008 382820
rect 234212 382780 234218 382792
rect 275002 382780 275008 382792
rect 275060 382780 275066 382832
rect 278958 382780 278964 382832
rect 279016 382820 279022 382832
rect 301682 382820 301688 382832
rect 279016 382792 301688 382820
rect 279016 382780 279022 382792
rect 301682 382780 301688 382792
rect 301740 382780 301746 382832
rect 234246 382712 234252 382764
rect 234304 382752 234310 382764
rect 280522 382752 280528 382764
rect 234304 382724 280528 382752
rect 234304 382712 234310 382724
rect 280522 382712 280528 382724
rect 280580 382712 280586 382764
rect 246114 382644 246120 382696
rect 246172 382684 246178 382696
rect 300762 382684 300768 382696
rect 246172 382656 300768 382684
rect 246172 382644 246178 382656
rect 300762 382644 300768 382656
rect 300820 382644 300826 382696
rect 174630 382576 174636 382628
rect 174688 382616 174694 382628
rect 258626 382616 258632 382628
rect 174688 382588 258632 382616
rect 174688 382576 174694 382588
rect 258626 382576 258632 382588
rect 258684 382576 258690 382628
rect 284478 382576 284484 382628
rect 284536 382616 284542 382628
rect 337378 382616 337384 382628
rect 284536 382588 337384 382616
rect 284536 382576 284542 382588
rect 337378 382576 337384 382588
rect 337436 382576 337442 382628
rect 94498 382508 94504 382560
rect 94556 382548 94562 382560
rect 267826 382548 267832 382560
rect 94556 382520 267832 382548
rect 94556 382508 94562 382520
rect 267826 382508 267832 382520
rect 267884 382508 267890 382560
rect 286134 382508 286140 382560
rect 286192 382548 286198 382560
rect 349246 382548 349252 382560
rect 286192 382520 349252 382548
rect 286192 382508 286198 382520
rect 349246 382508 349252 382520
rect 349304 382508 349310 382560
rect 91738 382440 91744 382492
rect 91796 382480 91802 382492
rect 266170 382480 266176 382492
rect 91796 382452 266176 382480
rect 91796 382440 91802 382452
rect 266170 382440 266176 382452
rect 266228 382440 266234 382492
rect 272518 382440 272524 382492
rect 272576 382480 272582 382492
rect 347866 382480 347872 382492
rect 272576 382452 347872 382480
rect 272576 382440 272582 382452
rect 347866 382440 347872 382452
rect 347924 382440 347930 382492
rect 233786 382372 233792 382424
rect 233844 382412 233850 382424
rect 265342 382412 265348 382424
rect 233844 382384 265348 382412
rect 233844 382372 233850 382384
rect 265342 382372 265348 382384
rect 265400 382372 265406 382424
rect 289078 382372 289084 382424
rect 289136 382412 289142 382424
rect 301590 382412 301596 382424
rect 289136 382384 301596 382412
rect 289136 382372 289142 382384
rect 301590 382372 301596 382384
rect 301648 382372 301654 382424
rect 235350 382304 235356 382356
rect 235408 382344 235414 382356
rect 265066 382344 265072 382356
rect 235408 382316 265072 382344
rect 235408 382304 235414 382316
rect 265066 382304 265072 382316
rect 265124 382304 265130 382356
rect 287238 382304 287244 382356
rect 287296 382344 287302 382356
rect 300302 382344 300308 382356
rect 287296 382316 300308 382344
rect 287296 382304 287302 382316
rect 300302 382304 300308 382316
rect 300360 382304 300366 382356
rect 232498 382236 232504 382288
rect 232556 382276 232562 382288
rect 265618 382276 265624 382288
rect 232556 382248 265624 382276
rect 232556 382236 232562 382248
rect 265618 382236 265624 382248
rect 265676 382236 265682 382288
rect 280062 382236 280068 382288
rect 280120 382276 280126 382288
rect 299474 382276 299480 382288
rect 280120 382248 299480 382276
rect 280120 382236 280126 382248
rect 299474 382236 299480 382248
rect 299532 382236 299538 382288
rect 257062 382004 257068 382016
rect 249766 381976 257068 382004
rect 242986 381896 242992 381948
rect 243044 381936 243050 381948
rect 248230 381936 248236 381948
rect 243044 381908 248236 381936
rect 243044 381896 243050 381908
rect 248230 381896 248236 381908
rect 248288 381896 248294 381948
rect 241606 381828 241612 381880
rect 241664 381868 241670 381880
rect 249766 381868 249794 381976
rect 257062 381964 257068 381976
rect 257120 381964 257126 382016
rect 263962 381964 263968 382016
rect 264020 382004 264026 382016
rect 265894 382004 265900 382016
rect 264020 381976 265900 382004
rect 264020 381964 264026 381976
rect 265894 381964 265900 381976
rect 265952 381964 265958 382016
rect 252922 381896 252928 381948
rect 252980 381936 252986 381948
rect 267274 381936 267280 381948
rect 252980 381908 267280 381936
rect 252980 381896 252986 381908
rect 267274 381896 267280 381908
rect 267332 381896 267338 381948
rect 268930 381868 268936 381880
rect 241664 381840 249794 381868
rect 260806 381840 268936 381868
rect 241664 381828 241670 381840
rect 245746 381760 245752 381812
rect 245804 381800 245810 381812
rect 256234 381800 256240 381812
rect 245804 381772 256240 381800
rect 245804 381760 245810 381772
rect 256234 381760 256240 381772
rect 256292 381760 256298 381812
rect 236822 381732 236828 381744
rect 234586 381704 236828 381732
rect 3694 381556 3700 381608
rect 3752 381596 3758 381608
rect 234586 381596 234614 381704
rect 236822 381692 236828 381704
rect 236880 381692 236886 381744
rect 243538 381692 243544 381744
rect 243596 381732 243602 381744
rect 247402 381732 247408 381744
rect 243596 381704 247408 381732
rect 243596 381692 243602 381704
rect 247402 381692 247408 381704
rect 247460 381692 247466 381744
rect 247678 381692 247684 381744
rect 247736 381732 247742 381744
rect 250714 381732 250720 381744
rect 247736 381704 250720 381732
rect 247736 381692 247742 381704
rect 250714 381692 250720 381704
rect 250772 381692 250778 381744
rect 255130 381692 255136 381744
rect 255188 381732 255194 381744
rect 259822 381732 259828 381744
rect 255188 381704 259828 381732
rect 255188 381692 255194 381704
rect 259822 381692 259828 381704
rect 259880 381692 259886 381744
rect 235902 381624 235908 381676
rect 235960 381664 235966 381676
rect 235960 381636 259454 381664
rect 235960 381624 235966 381636
rect 3752 381568 234614 381596
rect 3752 381556 3758 381568
rect 235534 381556 235540 381608
rect 235592 381596 235598 381608
rect 252922 381596 252928 381608
rect 235592 381568 252928 381596
rect 235592 381556 235598 381568
rect 252922 381556 252928 381568
rect 252980 381556 252986 381608
rect 3418 381488 3424 381540
rect 3476 381528 3482 381540
rect 239398 381528 239404 381540
rect 3476 381500 239404 381528
rect 3476 381488 3482 381500
rect 239398 381488 239404 381500
rect 239456 381488 239462 381540
rect 247678 381528 247684 381540
rect 241486 381500 247684 381528
rect 234430 381216 234436 381268
rect 234488 381256 234494 381268
rect 241486 381256 241514 381500
rect 247678 381488 247684 381500
rect 247736 381488 247742 381540
rect 250714 381488 250720 381540
rect 250772 381528 250778 381540
rect 259426 381528 259454 381636
rect 260806 381528 260834 381840
rect 268930 381828 268936 381840
rect 268988 381828 268994 381880
rect 264808 381772 273254 381800
rect 261202 381624 261208 381676
rect 261260 381664 261266 381676
rect 264808 381664 264836 381772
rect 270586 381732 270592 381744
rect 261260 381636 264836 381664
rect 270466 381704 270592 381732
rect 261260 381624 261266 381636
rect 270466 381596 270494 381704
rect 270586 381692 270592 381704
rect 270644 381692 270650 381744
rect 250772 381500 250852 381528
rect 259426 381500 260834 381528
rect 263888 381568 270494 381596
rect 250772 381488 250778 381500
rect 241606 381420 241612 381472
rect 241664 381420 241670 381472
rect 242986 381420 242992 381472
rect 243044 381420 243050 381472
rect 244366 381420 244372 381472
rect 244424 381420 244430 381472
rect 247402 381420 247408 381472
rect 247460 381460 247466 381472
rect 247460 381432 248184 381460
rect 247460 381420 247466 381432
rect 234488 381228 241514 381256
rect 234488 381216 234494 381228
rect 90450 381080 90456 381132
rect 90508 381120 90514 381132
rect 241624 381120 241652 381420
rect 90508 381092 241652 381120
rect 90508 381080 90514 381092
rect 3602 381012 3608 381064
rect 3660 381052 3666 381064
rect 3660 381024 234614 381052
rect 3660 381012 3666 381024
rect 234586 380916 234614 381024
rect 243004 380916 243032 381420
rect 244384 381188 244412 381420
rect 244384 381160 247356 381188
rect 234586 380888 243032 380916
rect 247328 380644 247356 381160
rect 248156 380780 248184 381432
rect 248230 381420 248236 381472
rect 248288 381420 248294 381472
rect 248248 381188 248276 381420
rect 250824 381256 250852 381500
rect 255130 381420 255136 381472
rect 255188 381420 255194 381472
rect 256234 381420 256240 381472
rect 256292 381420 256298 381472
rect 257062 381420 257068 381472
rect 257120 381460 257126 381472
rect 257120 381432 259454 381460
rect 257120 381420 257126 381432
rect 255148 381256 255176 381420
rect 250824 381228 255176 381256
rect 255424 381228 256188 381256
rect 248248 381160 251174 381188
rect 251146 381120 251174 381160
rect 255424 381120 255452 381228
rect 251146 381092 255452 381120
rect 256160 381052 256188 381228
rect 256252 381120 256280 381420
rect 259426 381256 259454 381432
rect 259822 381420 259828 381472
rect 259880 381420 259886 381472
rect 259840 381324 259868 381420
rect 263888 381324 263916 381568
rect 273226 381528 273254 381772
rect 275986 381704 285674 381732
rect 275986 381528 276014 381704
rect 276934 381624 276940 381676
rect 276992 381664 276998 381676
rect 282178 381664 282184 381676
rect 276992 381636 282184 381664
rect 276992 381624 276998 381636
rect 282178 381624 282184 381636
rect 282236 381624 282242 381676
rect 264808 381500 272104 381528
rect 273226 381500 276014 381528
rect 263962 381420 263968 381472
rect 264020 381420 264026 381472
rect 259840 381296 263916 381324
rect 263980 381256 264008 381420
rect 259426 381228 264008 381256
rect 264808 381120 264836 381500
rect 266722 381420 266728 381472
rect 266780 381420 266786 381472
rect 271966 381420 271972 381472
rect 272024 381420 272030 381472
rect 272076 381460 272104 381500
rect 277486 381488 277492 381540
rect 277544 381528 277550 381540
rect 285646 381528 285674 381704
rect 296806 381624 296812 381676
rect 296864 381664 296870 381676
rect 306374 381664 306380 381676
rect 296864 381636 306380 381664
rect 296864 381624 296870 381636
rect 306374 381624 306380 381636
rect 306432 381624 306438 381676
rect 293770 381556 293776 381608
rect 293828 381596 293834 381608
rect 579890 381596 579896 381608
rect 293828 381568 579896 381596
rect 293828 381556 293834 381568
rect 579890 381556 579896 381568
rect 579948 381556 579954 381608
rect 580074 381528 580080 381540
rect 277544 381500 281396 381528
rect 285646 381500 580080 381528
rect 277544 381488 277550 381500
rect 276934 381460 276940 381472
rect 272076 381432 276940 381460
rect 276934 381420 276940 381432
rect 276992 381420 276998 381472
rect 256252 381092 264836 381120
rect 266740 381052 266768 381420
rect 271984 381392 272012 381420
rect 271984 381364 275876 381392
rect 256160 381024 266768 381052
rect 275848 381052 275876 381364
rect 281368 381120 281396 381500
rect 580074 381488 580080 381500
rect 580132 381488 580138 381540
rect 282178 381420 282184 381472
rect 282236 381420 282242 381472
rect 283006 381420 283012 381472
rect 283064 381460 283070 381472
rect 283064 381432 287054 381460
rect 283064 381420 283070 381432
rect 282196 381392 282224 381420
rect 282196 381364 285674 381392
rect 285646 381188 285674 381364
rect 287026 381256 287054 381432
rect 300946 381256 300952 381268
rect 287026 381228 300952 381256
rect 300946 381216 300952 381228
rect 301004 381216 301010 381268
rect 301958 381188 301964 381200
rect 285646 381160 301964 381188
rect 301958 381148 301964 381160
rect 302016 381148 302022 381200
rect 300854 381120 300860 381132
rect 281368 381092 300860 381120
rect 300854 381080 300860 381092
rect 300912 381080 300918 381132
rect 344002 381052 344008 381064
rect 275848 381024 344008 381052
rect 344002 381012 344008 381024
rect 344060 381012 344066 381064
rect 580718 380984 580724 380996
rect 256068 380956 580724 380984
rect 256068 380780 256096 380956
rect 580718 380944 580724 380956
rect 580776 380944 580782 380996
rect 580902 380916 580908 380928
rect 248156 380752 256096 380780
rect 260806 380888 580908 380916
rect 260806 380644 260834 380888
rect 580902 380876 580908 380888
rect 580960 380876 580966 380928
rect 247328 380616 260834 380644
rect 300762 379448 300768 379500
rect 300820 379488 300826 379500
rect 580166 379488 580172 379500
rect 300820 379460 580172 379488
rect 300820 379448 300826 379460
rect 580166 379448 580172 379460
rect 580224 379448 580230 379500
rect 579982 378768 579988 378820
rect 580040 378808 580046 378820
rect 580810 378808 580816 378820
rect 580040 378780 580816 378808
rect 580040 378768 580046 378780
rect 580810 378768 580816 378780
rect 580868 378768 580874 378820
rect 3142 372512 3148 372564
rect 3200 372552 3206 372564
rect 174630 372552 174636 372564
rect 3200 372524 174636 372552
rect 3200 372512 3206 372524
rect 174630 372512 174636 372524
rect 174688 372512 174694 372564
rect 301958 353200 301964 353252
rect 302016 353240 302022 353252
rect 579982 353240 579988 353252
rect 302016 353212 579988 353240
rect 302016 353200 302022 353212
rect 579982 353200 579988 353212
rect 580040 353200 580046 353252
rect 2958 346332 2964 346384
rect 3016 346372 3022 346384
rect 235166 346372 235172 346384
rect 3016 346344 235172 346372
rect 3016 346332 3022 346344
rect 235166 346332 235172 346344
rect 235224 346332 235230 346384
rect 244090 338512 244096 338564
rect 244148 338552 244154 338564
rect 244148 338524 251174 338552
rect 244148 338512 244154 338524
rect 251146 338348 251174 338524
rect 251146 338320 256418 338348
rect 244734 338036 244740 338088
rect 244792 338076 244798 338088
rect 244792 338048 249886 338076
rect 244792 338036 244798 338048
rect 242986 337968 242992 338020
rect 243044 338008 243050 338020
rect 243044 337980 247310 338008
rect 243044 337968 243050 337980
rect 244458 337900 244464 337952
rect 244516 337940 244522 337952
rect 245608 337940 245614 337952
rect 244516 337912 245614 337940
rect 244516 337900 244522 337912
rect 245608 337900 245614 337912
rect 245666 337900 245672 337952
rect 245700 337900 245706 337952
rect 245758 337900 245764 337952
rect 245884 337900 245890 337952
rect 245942 337900 245948 337952
rect 246252 337900 246258 337952
rect 246310 337900 246316 337952
rect 246436 337900 246442 337952
rect 246494 337900 246500 337952
rect 246712 337900 246718 337952
rect 246770 337900 246776 337952
rect 246804 337900 246810 337952
rect 246862 337900 246868 337952
rect 246896 337900 246902 337952
rect 246954 337900 246960 337952
rect 247080 337900 247086 337952
rect 247138 337900 247144 337952
rect 247172 337900 247178 337952
rect 247230 337900 247236 337952
rect 247282 337940 247310 337980
rect 247466 337980 248782 338008
rect 247356 337940 247362 337952
rect 247282 337912 247362 337940
rect 247356 337900 247362 337912
rect 247414 337900 247420 337952
rect 245102 337832 245108 337884
rect 245160 337872 245166 337884
rect 245718 337872 245746 337900
rect 245160 337844 245746 337872
rect 245160 337832 245166 337844
rect 244274 337764 244280 337816
rect 244332 337804 244338 337816
rect 245516 337804 245522 337816
rect 244332 337776 245522 337804
rect 244332 337764 244338 337776
rect 245516 337764 245522 337776
rect 245574 337764 245580 337816
rect 245902 337748 245930 337900
rect 245902 337708 245936 337748
rect 245930 337696 245936 337708
rect 245988 337696 245994 337748
rect 246022 337628 246028 337680
rect 246080 337668 246086 337680
rect 246270 337668 246298 337900
rect 246080 337640 246298 337668
rect 246080 337628 246086 337640
rect 246454 337544 246482 337900
rect 246620 337872 246626 337884
rect 246592 337832 246626 337872
rect 246678 337832 246684 337884
rect 246592 337612 246620 337832
rect 246730 337804 246758 337900
rect 246684 337776 246758 337804
rect 246684 337748 246712 337776
rect 246822 337748 246850 337900
rect 246666 337696 246672 337748
rect 246724 337696 246730 337748
rect 246758 337696 246764 337748
rect 246816 337708 246850 337748
rect 246816 337696 246822 337708
rect 246574 337560 246580 337612
rect 246632 337560 246638 337612
rect 246454 337504 246488 337544
rect 246482 337492 246488 337504
rect 246540 337492 246546 337544
rect 245010 337424 245016 337476
rect 245068 337464 245074 337476
rect 246914 337464 246942 337900
rect 247098 337872 247126 337900
rect 247052 337844 247126 337872
rect 247052 337736 247080 337844
rect 247190 337816 247218 337900
rect 247264 337832 247270 337884
rect 247322 337872 247328 337884
rect 247466 337872 247494 337980
rect 248754 337952 248782 337980
rect 249858 337952 249886 338048
rect 254918 337980 255544 338008
rect 254918 337952 254946 337980
rect 247816 337900 247822 337952
rect 247874 337940 247880 337952
rect 248276 337940 248282 337952
rect 247874 337900 247908 337940
rect 247322 337832 247356 337872
rect 247126 337764 247132 337816
rect 247184 337776 247218 337816
rect 247184 337764 247190 337776
rect 247328 337748 247356 337832
rect 247420 337844 247494 337872
rect 247420 337816 247448 337844
rect 247632 337832 247638 337884
rect 247690 337832 247696 337884
rect 247402 337764 247408 337816
rect 247460 337764 247466 337816
rect 247650 337804 247678 337832
rect 247880 337816 247908 337900
rect 248248 337900 248282 337940
rect 248334 337900 248340 337952
rect 248368 337900 248374 337952
rect 248426 337900 248432 337952
rect 248644 337940 248650 337952
rect 248616 337900 248650 337940
rect 248702 337900 248708 337952
rect 248736 337900 248742 337952
rect 248794 337900 248800 337952
rect 248828 337900 248834 337952
rect 248886 337900 248892 337952
rect 248920 337900 248926 337952
rect 248978 337900 248984 337952
rect 249104 337940 249110 337952
rect 249076 337900 249110 337940
rect 249162 337900 249168 337952
rect 249196 337900 249202 337952
rect 249254 337900 249260 337952
rect 249288 337900 249294 337952
rect 249346 337940 249352 337952
rect 249656 337940 249662 337952
rect 249346 337900 249380 337940
rect 248000 337832 248006 337884
rect 248058 337832 248064 337884
rect 248092 337832 248098 337884
rect 248150 337832 248156 337884
rect 247512 337776 247678 337804
rect 247218 337736 247224 337748
rect 247052 337708 247224 337736
rect 247218 337696 247224 337708
rect 247276 337696 247282 337748
rect 247310 337696 247316 337748
rect 247368 337696 247374 337748
rect 247218 337560 247224 337612
rect 247276 337600 247282 337612
rect 247512 337600 247540 337776
rect 247862 337764 247868 337816
rect 247920 337764 247926 337816
rect 248018 337736 248046 337832
rect 247604 337708 248046 337736
rect 247604 337680 247632 337708
rect 247586 337628 247592 337680
rect 247644 337628 247650 337680
rect 248110 337668 248138 337832
rect 247788 337640 248138 337668
rect 247788 337612 247816 337640
rect 247276 337572 247540 337600
rect 247276 337560 247282 337572
rect 247770 337560 247776 337612
rect 247828 337560 247834 337612
rect 248248 337544 248276 337900
rect 248386 337680 248414 337900
rect 248460 337832 248466 337884
rect 248518 337872 248524 337884
rect 248518 337832 248552 337872
rect 248524 337748 248552 337832
rect 248506 337696 248512 337748
rect 248564 337696 248570 337748
rect 248616 337680 248644 337900
rect 248846 337816 248874 337900
rect 248782 337764 248788 337816
rect 248840 337776 248874 337816
rect 248840 337764 248846 337776
rect 248938 337748 248966 337900
rect 248874 337696 248880 337748
rect 248932 337708 248966 337748
rect 248932 337696 248938 337708
rect 248322 337628 248328 337680
rect 248380 337640 248414 337680
rect 248380 337628 248386 337640
rect 248598 337628 248604 337680
rect 248656 337628 248662 337680
rect 249076 337600 249104 337900
rect 249214 337680 249242 337900
rect 249150 337628 249156 337680
rect 249208 337640 249242 337680
rect 249208 337628 249214 337640
rect 249242 337600 249248 337612
rect 249076 337572 249248 337600
rect 249242 337560 249248 337572
rect 249300 337560 249306 337612
rect 249352 337544 249380 337900
rect 249628 337900 249662 337940
rect 249714 337900 249720 337952
rect 249748 337900 249754 337952
rect 249806 337900 249812 337952
rect 249840 337900 249846 337952
rect 249898 337900 249904 337952
rect 250024 337900 250030 337952
rect 250082 337900 250088 337952
rect 250116 337900 250122 337952
rect 250174 337900 250180 337952
rect 250208 337900 250214 337952
rect 250266 337900 250272 337952
rect 250760 337900 250766 337952
rect 250818 337900 250824 337952
rect 250852 337900 250858 337952
rect 250910 337900 250916 337952
rect 251036 337900 251042 337952
rect 251094 337900 251100 337952
rect 251404 337900 251410 337952
rect 251462 337900 251468 337952
rect 251680 337900 251686 337952
rect 251738 337900 251744 337952
rect 252048 337900 252054 337952
rect 252106 337900 252112 337952
rect 252324 337900 252330 337952
rect 252382 337940 252388 337952
rect 253428 337940 253434 337952
rect 252382 337900 252416 337940
rect 249472 337804 249478 337816
rect 249444 337764 249478 337804
rect 249530 337764 249536 337816
rect 248230 337492 248236 337544
rect 248288 337492 248294 337544
rect 249334 337492 249340 337544
rect 249392 337492 249398 337544
rect 245068 337436 246942 337464
rect 245068 337424 245074 337436
rect 248138 337424 248144 337476
rect 248196 337464 248202 337476
rect 249444 337464 249472 337764
rect 249628 337748 249656 337900
rect 249766 337872 249794 337900
rect 249720 337844 249794 337872
rect 249610 337696 249616 337748
rect 249668 337696 249674 337748
rect 249720 337680 249748 337844
rect 250042 337816 250070 337900
rect 249978 337764 249984 337816
rect 250036 337776 250070 337816
rect 250036 337764 250042 337776
rect 249702 337628 249708 337680
rect 249760 337628 249766 337680
rect 249518 337560 249524 337612
rect 249576 337600 249582 337612
rect 250134 337600 250162 337900
rect 250226 337816 250254 337900
rect 250576 337832 250582 337884
rect 250634 337832 250640 337884
rect 250208 337764 250214 337816
rect 250266 337764 250272 337816
rect 250594 337612 250622 337832
rect 250778 337612 250806 337900
rect 249576 337572 250162 337600
rect 249576 337560 249582 337572
rect 250530 337560 250536 337612
rect 250588 337572 250622 337612
rect 250588 337560 250594 337572
rect 250714 337560 250720 337612
rect 250772 337572 250806 337612
rect 250772 337560 250778 337572
rect 249886 337492 249892 337544
rect 249944 337532 249950 337544
rect 250870 337532 250898 337900
rect 251054 337680 251082 337900
rect 251128 337832 251134 337884
rect 251186 337872 251192 337884
rect 251312 337872 251318 337884
rect 251186 337832 251220 337872
rect 251192 337748 251220 337832
rect 251284 337832 251318 337872
rect 251370 337832 251376 337884
rect 251174 337696 251180 337748
rect 251232 337696 251238 337748
rect 250990 337628 250996 337680
rect 251048 337640 251082 337680
rect 251048 337628 251054 337640
rect 251082 337560 251088 337612
rect 251140 337600 251146 337612
rect 251284 337600 251312 337832
rect 251422 337612 251450 337900
rect 251698 337816 251726 337900
rect 251864 337832 251870 337884
rect 251922 337832 251928 337884
rect 251634 337764 251640 337816
rect 251692 337776 251726 337816
rect 251692 337764 251698 337776
rect 251882 337736 251910 337832
rect 252066 337816 252094 337900
rect 252232 337832 252238 337884
rect 252290 337832 252296 337884
rect 252002 337764 252008 337816
rect 252060 337776 252094 337816
rect 252060 337764 252066 337776
rect 251560 337708 251910 337736
rect 251560 337612 251588 337708
rect 251140 337572 251312 337600
rect 251140 337560 251146 337572
rect 251358 337560 251364 337612
rect 251416 337572 251450 337612
rect 251416 337560 251422 337572
rect 251542 337560 251548 337612
rect 251600 337560 251606 337612
rect 251726 337560 251732 337612
rect 251784 337600 251790 337612
rect 252250 337600 252278 337832
rect 252388 337680 252416 337900
rect 252802 337912 253434 337940
rect 252600 337872 252606 337884
rect 252480 337844 252606 337872
rect 252370 337628 252376 337680
rect 252428 337628 252434 337680
rect 251784 337572 252278 337600
rect 251784 337560 251790 337572
rect 249944 337504 250898 337532
rect 249944 337492 249950 337504
rect 251450 337492 251456 337544
rect 251508 337532 251514 337544
rect 252480 337532 252508 337844
rect 252600 337832 252606 337844
rect 252658 337832 252664 337884
rect 252802 337736 252830 337912
rect 253428 337900 253434 337912
rect 253486 337900 253492 337952
rect 253888 337900 253894 337952
rect 253946 337900 253952 337952
rect 254900 337900 254906 337952
rect 254958 337900 254964 337952
rect 255084 337900 255090 337952
rect 255142 337900 255148 337952
rect 255176 337900 255182 337952
rect 255234 337900 255240 337952
rect 255268 337900 255274 337952
rect 255326 337900 255332 337952
rect 255360 337900 255366 337952
rect 255418 337900 255424 337952
rect 253152 337832 253158 337884
rect 253210 337832 253216 337884
rect 253244 337832 253250 337884
rect 253302 337832 253308 337884
rect 253612 337832 253618 337884
rect 253670 337832 253676 337884
rect 253170 337804 253198 337832
rect 252572 337708 252830 337736
rect 252894 337776 253198 337804
rect 252572 337612 252600 337708
rect 252894 337612 252922 337776
rect 253262 337736 253290 337832
rect 253124 337708 253290 337736
rect 253124 337680 253152 337708
rect 253106 337628 253112 337680
rect 253164 337628 253170 337680
rect 253290 337628 253296 337680
rect 253348 337668 253354 337680
rect 253630 337668 253658 337832
rect 253906 337748 253934 337900
rect 254256 337872 254262 337884
rect 254228 337832 254262 337872
rect 254314 337832 254320 337884
rect 254440 337832 254446 337884
rect 254498 337832 254504 337884
rect 255102 337872 255130 337900
rect 255056 337844 255130 337872
rect 254072 337764 254078 337816
rect 254130 337764 254136 337816
rect 253906 337708 253940 337748
rect 253934 337696 253940 337708
rect 253992 337696 253998 337748
rect 253348 337640 253658 337668
rect 254090 337680 254118 337764
rect 254228 337748 254256 337832
rect 254210 337696 254216 337748
rect 254268 337696 254274 337748
rect 254090 337640 254124 337680
rect 253348 337628 253354 337640
rect 254118 337628 254124 337640
rect 254176 337628 254182 337680
rect 254458 337668 254486 337832
rect 255056 337816 255084 337844
rect 255194 337816 255222 337900
rect 254532 337764 254538 337816
rect 254590 337764 254596 337816
rect 254624 337764 254630 337816
rect 254682 337764 254688 337816
rect 254716 337764 254722 337816
rect 254774 337764 254780 337816
rect 255038 337764 255044 337816
rect 255096 337764 255102 337816
rect 255130 337764 255136 337816
rect 255188 337776 255222 337816
rect 255188 337764 255194 337776
rect 254320 337640 254486 337668
rect 254320 337612 254348 337640
rect 252554 337560 252560 337612
rect 252612 337560 252618 337612
rect 252830 337560 252836 337612
rect 252888 337572 252922 337612
rect 252888 337560 252894 337572
rect 254302 337560 254308 337612
rect 254360 337560 254366 337612
rect 254550 337600 254578 337764
rect 254504 337572 254578 337600
rect 254642 337612 254670 337764
rect 254734 337680 254762 337764
rect 255286 337748 255314 337900
rect 255222 337696 255228 337748
rect 255280 337708 255314 337748
rect 255280 337696 255286 337708
rect 254734 337640 254768 337680
rect 254762 337628 254768 337640
rect 254820 337628 254826 337680
rect 255378 337612 255406 337900
rect 255516 337680 255544 337980
rect 256188 337900 256194 337952
rect 256246 337900 256252 337952
rect 255498 337628 255504 337680
rect 255556 337628 255562 337680
rect 254642 337572 254676 337612
rect 254504 337544 254532 337572
rect 254670 337560 254676 337572
rect 254728 337560 254734 337612
rect 255314 337560 255320 337612
rect 255372 337572 255406 337612
rect 255372 337560 255378 337572
rect 251508 337504 252508 337532
rect 251508 337492 251514 337504
rect 254486 337492 254492 337544
rect 254544 337492 254550 337544
rect 256206 337532 256234 337900
rect 256390 337600 256418 338320
rect 288406 338320 292574 338348
rect 288406 338280 288434 338320
rect 280126 338252 288434 338280
rect 292546 338280 292574 338320
rect 430574 338280 430580 338292
rect 292546 338252 430580 338280
rect 274606 338184 275784 338212
rect 274606 338076 274634 338184
rect 270282 338048 274634 338076
rect 270282 337952 270310 338048
rect 273778 337980 274634 338008
rect 273778 337952 273806 337980
rect 257292 337900 257298 337952
rect 257350 337900 257356 337952
rect 257384 337900 257390 337952
rect 257442 337900 257448 337952
rect 257568 337900 257574 337952
rect 257626 337900 257632 337952
rect 257936 337900 257942 337952
rect 257994 337900 258000 337952
rect 258396 337940 258402 337952
rect 258276 337912 258402 337940
rect 256648 337872 256654 337884
rect 256528 337844 256654 337872
rect 256390 337572 256464 337600
rect 256436 337544 256464 337572
rect 254596 337504 256234 337532
rect 248196 337436 249472 337464
rect 248196 337424 248202 337436
rect 250346 337424 250352 337476
rect 250404 337464 250410 337476
rect 250898 337464 250904 337476
rect 250404 337436 250904 337464
rect 250404 337424 250410 337436
rect 250898 337424 250904 337436
rect 250956 337424 250962 337476
rect 254596 337464 254624 337504
rect 256418 337492 256424 337544
rect 256476 337492 256482 337544
rect 253998 337436 254624 337464
rect 139394 337356 139400 337408
rect 139452 337396 139458 337408
rect 253998 337396 254026 337436
rect 255682 337424 255688 337476
rect 255740 337464 255746 337476
rect 256528 337464 256556 337844
rect 256648 337832 256654 337844
rect 256706 337832 256712 337884
rect 256832 337872 256838 337884
rect 256758 337844 256838 337872
rect 256758 337804 256786 337844
rect 256832 337832 256838 337844
rect 256890 337832 256896 337884
rect 256712 337776 256786 337804
rect 256712 337600 256740 337776
rect 257310 337736 257338 337900
rect 256988 337708 257338 337736
rect 257402 337748 257430 337900
rect 257402 337708 257436 337748
rect 256786 337600 256792 337612
rect 256712 337572 256792 337600
rect 256786 337560 256792 337572
rect 256844 337560 256850 337612
rect 256988 337476 257016 337708
rect 257430 337696 257436 337708
rect 257488 337696 257494 337748
rect 257338 337560 257344 337612
rect 257396 337600 257402 337612
rect 257586 337600 257614 337900
rect 257660 337832 257666 337884
rect 257718 337832 257724 337884
rect 257396 337572 257614 337600
rect 257396 337560 257402 337572
rect 255740 337436 256556 337464
rect 255740 337424 255746 337436
rect 256970 337424 256976 337476
rect 257028 337424 257034 337476
rect 139452 337368 244964 337396
rect 139452 337356 139458 337368
rect 81434 337288 81440 337340
rect 81492 337328 81498 337340
rect 244936 337328 244964 337368
rect 246500 337368 254026 337396
rect 246500 337328 246528 337368
rect 256878 337356 256884 337408
rect 256936 337396 256942 337408
rect 257678 337396 257706 337832
rect 257844 337764 257850 337816
rect 257902 337764 257908 337816
rect 257862 337680 257890 337764
rect 257798 337628 257804 337680
rect 257856 337640 257890 337680
rect 257856 337628 257862 337640
rect 257954 337612 257982 337900
rect 258120 337764 258126 337816
rect 258178 337764 258184 337816
rect 258138 337680 258166 337764
rect 258074 337628 258080 337680
rect 258132 337640 258166 337680
rect 258132 337628 258138 337640
rect 257890 337560 257896 337612
rect 257948 337572 257982 337612
rect 257948 337560 257954 337572
rect 258276 337544 258304 337912
rect 258396 337900 258402 337912
rect 258454 337900 258460 337952
rect 258488 337900 258494 337952
rect 258546 337900 258552 337952
rect 258672 337900 258678 337952
rect 258730 337900 258736 337952
rect 258856 337900 258862 337952
rect 258914 337900 258920 337952
rect 258948 337900 258954 337952
rect 259006 337900 259012 337952
rect 259224 337900 259230 337952
rect 259282 337900 259288 337952
rect 259408 337900 259414 337952
rect 259466 337900 259472 337952
rect 259500 337900 259506 337952
rect 259558 337900 259564 337952
rect 259592 337900 259598 337952
rect 259650 337900 259656 337952
rect 259868 337900 259874 337952
rect 259926 337900 259932 337952
rect 259960 337900 259966 337952
rect 260018 337900 260024 337952
rect 260236 337900 260242 337952
rect 260294 337900 260300 337952
rect 260420 337900 260426 337952
rect 260478 337900 260484 337952
rect 260512 337900 260518 337952
rect 260570 337900 260576 337952
rect 261248 337900 261254 337952
rect 261306 337940 261312 337952
rect 261306 337900 261340 337940
rect 261616 337900 261622 337952
rect 261674 337900 261680 337952
rect 261708 337900 261714 337952
rect 261766 337900 261772 337952
rect 262076 337940 262082 337952
rect 262048 337900 262082 337940
rect 262134 337900 262140 337952
rect 262260 337900 262266 337952
rect 262318 337900 262324 337952
rect 262720 337900 262726 337952
rect 262778 337900 262784 337952
rect 262904 337940 262910 337952
rect 262830 337912 262910 337940
rect 258506 337872 258534 337900
rect 258368 337844 258534 337872
rect 258368 337680 258396 337844
rect 258442 337764 258448 337816
rect 258500 337804 258506 337816
rect 258690 337804 258718 337900
rect 258500 337776 258718 337804
rect 258500 337764 258506 337776
rect 258350 337628 258356 337680
rect 258408 337628 258414 337680
rect 258874 337612 258902 337900
rect 258810 337560 258816 337612
rect 258868 337572 258902 337612
rect 258966 337612 258994 337900
rect 258966 337572 259000 337612
rect 258868 337560 258874 337572
rect 258994 337560 259000 337572
rect 259052 337560 259058 337612
rect 258258 337492 258264 337544
rect 258316 337492 258322 337544
rect 258534 337492 258540 337544
rect 258592 337532 258598 337544
rect 259242 337532 259270 337900
rect 259426 337872 259454 337900
rect 259380 337844 259454 337872
rect 259380 337680 259408 337844
rect 259518 337816 259546 337900
rect 259454 337764 259460 337816
rect 259512 337776 259546 337816
rect 259512 337764 259518 337776
rect 259610 337748 259638 337900
rect 259684 337832 259690 337884
rect 259742 337832 259748 337884
rect 259546 337696 259552 337748
rect 259604 337708 259638 337748
rect 259604 337696 259610 337708
rect 259362 337628 259368 337680
rect 259420 337628 259426 337680
rect 259702 337668 259730 337832
rect 259886 337816 259914 337900
rect 259978 337872 260006 337900
rect 259978 337844 260144 337872
rect 259868 337764 259874 337816
rect 259926 337764 259932 337816
rect 259702 337640 259960 337668
rect 258592 337504 259270 337532
rect 258592 337492 258598 337504
rect 259638 337492 259644 337544
rect 259696 337532 259702 337544
rect 259932 337532 259960 337640
rect 259696 337504 259960 337532
rect 259696 337492 259702 337504
rect 259822 337424 259828 337476
rect 259880 337464 259886 337476
rect 260116 337464 260144 337844
rect 260254 337680 260282 337900
rect 260190 337628 260196 337680
rect 260248 337640 260282 337680
rect 260248 337628 260254 337640
rect 259880 337436 260144 337464
rect 260438 337476 260466 337900
rect 260530 337544 260558 337900
rect 261156 337832 261162 337884
rect 261214 337872 261220 337884
rect 261214 337832 261248 337872
rect 260696 337764 260702 337816
rect 260754 337764 260760 337816
rect 260530 337504 260564 337544
rect 260558 337492 260564 337504
rect 260616 337492 260622 337544
rect 260714 337476 260742 337764
rect 261220 337748 261248 337832
rect 261202 337696 261208 337748
rect 261260 337696 261266 337748
rect 261110 337560 261116 337612
rect 261168 337600 261174 337612
rect 261312 337600 261340 337900
rect 261634 337736 261662 337900
rect 261168 337572 261340 337600
rect 261588 337708 261662 337736
rect 261588 337600 261616 337708
rect 261726 337680 261754 337900
rect 262048 337816 262076 337900
rect 262168 337872 262174 337884
rect 262140 337832 262174 337872
rect 262226 337832 262232 337884
rect 262030 337764 262036 337816
rect 262088 337764 262094 337816
rect 261662 337628 261668 337680
rect 261720 337640 261754 337680
rect 261720 337628 261726 337640
rect 261938 337600 261944 337612
rect 261588 337572 261944 337600
rect 261168 337560 261174 337572
rect 261938 337560 261944 337572
rect 261996 337560 262002 337612
rect 261202 337492 261208 337544
rect 261260 337532 261266 337544
rect 262140 337532 262168 337832
rect 262278 337748 262306 337900
rect 262444 337764 262450 337816
rect 262502 337764 262508 337816
rect 262214 337696 262220 337748
rect 262272 337708 262306 337748
rect 262272 337696 262278 337708
rect 262462 337600 262490 337764
rect 262582 337600 262588 337612
rect 262462 337572 262588 337600
rect 262582 337560 262588 337572
rect 262640 337560 262646 337612
rect 261260 337504 262168 337532
rect 261260 337492 261266 337504
rect 262490 337492 262496 337544
rect 262548 337532 262554 337544
rect 262738 337532 262766 337900
rect 262548 337504 262766 337532
rect 262548 337492 262554 337504
rect 260438 337436 260472 337476
rect 259880 337424 259886 337436
rect 260466 337424 260472 337436
rect 260524 337424 260530 337476
rect 260650 337424 260656 337476
rect 260708 337436 260742 337476
rect 260708 337424 260714 337436
rect 256936 337368 257706 337396
rect 256936 337356 256942 337368
rect 259914 337356 259920 337408
rect 259972 337396 259978 337408
rect 262830 337396 262858 337912
rect 262904 337900 262910 337912
rect 262962 337900 262968 337952
rect 262996 337900 263002 337952
rect 263054 337900 263060 337952
rect 263088 337900 263094 337952
rect 263146 337900 263152 337952
rect 263548 337900 263554 337952
rect 263606 337900 263612 337952
rect 263640 337900 263646 337952
rect 263698 337900 263704 337952
rect 264008 337900 264014 337952
rect 264066 337900 264072 337952
rect 265480 337900 265486 337952
rect 265538 337900 265544 337952
rect 266952 337940 266958 337952
rect 265820 337912 266958 337940
rect 263014 337816 263042 337900
rect 262950 337764 262956 337816
rect 263008 337776 263042 337816
rect 263008 337764 263014 337776
rect 263106 337736 263134 337900
rect 263272 337764 263278 337816
rect 263330 337764 263336 337816
rect 263106 337708 263180 337736
rect 263152 337680 263180 337708
rect 263134 337628 263140 337680
rect 263192 337628 263198 337680
rect 263290 337476 263318 337764
rect 263566 337476 263594 337900
rect 263226 337424 263232 337476
rect 263284 337436 263318 337476
rect 263284 337424 263290 337436
rect 263502 337424 263508 337476
rect 263560 337436 263594 337476
rect 263658 337476 263686 337900
rect 263824 337832 263830 337884
rect 263882 337832 263888 337884
rect 263842 337748 263870 337832
rect 263842 337708 263876 337748
rect 263870 337696 263876 337708
rect 263928 337696 263934 337748
rect 264026 337680 264054 337900
rect 264652 337832 264658 337884
rect 264710 337832 264716 337884
rect 264744 337832 264750 337884
rect 264802 337832 264808 337884
rect 265020 337832 265026 337884
rect 265078 337872 265084 337884
rect 265078 337832 265112 337872
rect 265296 337832 265302 337884
rect 265354 337872 265360 337884
rect 265354 337832 265388 337872
rect 264192 337764 264198 337816
rect 264250 337764 264256 337816
rect 264376 337764 264382 337816
rect 264434 337764 264440 337816
rect 264026 337640 264060 337680
rect 264054 337628 264060 337640
rect 264112 337628 264118 337680
rect 264210 337668 264238 337764
rect 264394 337680 264422 337764
rect 264210 337640 264284 337668
rect 264394 337640 264428 337680
rect 263658 337436 263692 337476
rect 263560 337424 263566 337436
rect 263686 337424 263692 337436
rect 263744 337424 263750 337476
rect 264256 337408 264284 337640
rect 264422 337628 264428 337640
rect 264480 337628 264486 337680
rect 264670 337600 264698 337832
rect 264348 337572 264698 337600
rect 259972 337368 262858 337396
rect 259972 337356 259978 337368
rect 264238 337356 264244 337408
rect 264296 337356 264302 337408
rect 81492 337300 244274 337328
rect 244936 337300 246528 337328
rect 81492 337288 81498 337300
rect 26234 337220 26240 337272
rect 26292 337260 26298 337272
rect 242986 337260 242992 337272
rect 26292 337232 242992 337260
rect 26292 337220 26298 337232
rect 242986 337220 242992 337232
rect 243044 337220 243050 337272
rect 244246 337260 244274 337300
rect 248966 337288 248972 337340
rect 249024 337328 249030 337340
rect 253934 337328 253940 337340
rect 249024 337300 253940 337328
rect 249024 337288 249030 337300
rect 253934 337288 253940 337300
rect 253992 337288 253998 337340
rect 264146 337288 264152 337340
rect 264204 337328 264210 337340
rect 264348 337328 264376 337572
rect 264606 337492 264612 337544
rect 264664 337532 264670 337544
rect 264762 337532 264790 337832
rect 265084 337748 265112 337832
rect 265360 337748 265388 337832
rect 265066 337696 265072 337748
rect 265124 337696 265130 337748
rect 265342 337696 265348 337748
rect 265400 337696 265406 337748
rect 264664 337504 264790 337532
rect 264664 337492 264670 337504
rect 265158 337492 265164 337544
rect 265216 337532 265222 337544
rect 265498 337532 265526 337900
rect 265664 337872 265670 337884
rect 265636 337832 265670 337872
rect 265722 337832 265728 337884
rect 265636 337680 265664 337832
rect 265710 337696 265716 337748
rect 265768 337696 265774 337748
rect 265618 337628 265624 337680
rect 265676 337628 265682 337680
rect 265728 337612 265756 337696
rect 265710 337560 265716 337612
rect 265768 337560 265774 337612
rect 265216 337504 265526 337532
rect 265216 337492 265222 337504
rect 264974 337424 264980 337476
rect 265032 337464 265038 337476
rect 265820 337464 265848 337912
rect 266952 337900 266958 337912
rect 267010 337900 267016 337952
rect 267044 337900 267050 337952
rect 267102 337900 267108 337952
rect 267136 337900 267142 337952
rect 267194 337900 267200 337952
rect 267504 337900 267510 337952
rect 267562 337900 267568 337952
rect 268056 337900 268062 337952
rect 268114 337900 268120 337952
rect 269068 337900 269074 337952
rect 269126 337900 269132 337952
rect 269344 337900 269350 337952
rect 269402 337900 269408 337952
rect 269712 337900 269718 337952
rect 269770 337900 269776 337952
rect 269804 337900 269810 337952
rect 269862 337940 269868 337952
rect 269862 337912 270218 337940
rect 269862 337900 269868 337912
rect 265940 337832 265946 337884
rect 265998 337832 266004 337884
rect 266492 337832 266498 337884
rect 266550 337832 266556 337884
rect 266584 337832 266590 337884
rect 266642 337832 266648 337884
rect 265958 337476 265986 337832
rect 266078 337560 266084 337612
rect 266136 337560 266142 337612
rect 265032 337436 265848 337464
rect 265032 337424 265038 337436
rect 265894 337424 265900 337476
rect 265952 337436 265986 337476
rect 265952 337424 265958 337436
rect 265802 337356 265808 337408
rect 265860 337396 265866 337408
rect 266096 337396 266124 337560
rect 266510 337532 266538 337832
rect 266602 337748 266630 337832
rect 267062 337816 267090 337900
rect 266998 337764 267004 337816
rect 267056 337776 267090 337816
rect 267056 337764 267062 337776
rect 267154 337748 267182 337900
rect 267228 337832 267234 337884
rect 267286 337832 267292 337884
rect 267320 337832 267326 337884
rect 267378 337832 267384 337884
rect 266602 337708 266636 337748
rect 266630 337696 266636 337708
rect 266688 337696 266694 337748
rect 267090 337696 267096 337748
rect 267148 337708 267182 337748
rect 267148 337696 267154 337708
rect 267246 337680 267274 337832
rect 267182 337628 267188 337680
rect 267240 337640 267274 337680
rect 267240 337628 267246 337640
rect 267338 337612 267366 337832
rect 267522 337680 267550 337900
rect 267458 337628 267464 337680
rect 267516 337640 267550 337680
rect 267516 337628 267522 337640
rect 267338 337572 267372 337612
rect 267366 337560 267372 337572
rect 267424 337560 267430 337612
rect 268074 337600 268102 337900
rect 268332 337832 268338 337884
rect 268390 337832 268396 337884
rect 268792 337832 268798 337884
rect 268850 337832 268856 337884
rect 267752 337572 268102 337600
rect 268350 337600 268378 337832
rect 268350 337572 268516 337600
rect 267752 337544 267780 337572
rect 268488 337544 268516 337572
rect 266630 337532 266636 337544
rect 266510 337504 266636 337532
rect 266630 337492 266636 337504
rect 266688 337492 266694 337544
rect 267734 337492 267740 337544
rect 267792 337492 267798 337544
rect 268470 337492 268476 337544
rect 268528 337492 268534 337544
rect 268102 337424 268108 337476
rect 268160 337464 268166 337476
rect 268810 337464 268838 337832
rect 268930 337628 268936 337680
rect 268988 337668 268994 337680
rect 269086 337668 269114 337900
rect 269160 337832 269166 337884
rect 269218 337832 269224 337884
rect 268988 337640 269114 337668
rect 268988 337628 268994 337640
rect 269178 337544 269206 337832
rect 269362 337680 269390 337900
rect 269730 337872 269758 337900
rect 269298 337628 269304 337680
rect 269356 337640 269390 337680
rect 269454 337844 269758 337872
rect 269454 337680 269482 337844
rect 270080 337832 270086 337884
rect 270138 337832 270144 337884
rect 269528 337764 269534 337816
rect 269586 337804 269592 337816
rect 269758 337804 269764 337816
rect 269586 337776 269764 337804
rect 269586 337764 269592 337776
rect 269758 337764 269764 337776
rect 269816 337764 269822 337816
rect 269454 337640 269488 337680
rect 269356 337628 269362 337640
rect 269482 337628 269488 337640
rect 269540 337628 269546 337680
rect 269574 337628 269580 337680
rect 269632 337668 269638 337680
rect 270098 337668 270126 337832
rect 269632 337640 270126 337668
rect 269632 337628 269638 337640
rect 270034 337560 270040 337612
rect 270092 337600 270098 337612
rect 270190 337600 270218 337912
rect 270264 337900 270270 337952
rect 270322 337900 270328 337952
rect 270356 337900 270362 337952
rect 270414 337900 270420 337952
rect 270724 337900 270730 337952
rect 270782 337900 270788 337952
rect 271092 337900 271098 337952
rect 271150 337900 271156 337952
rect 271184 337900 271190 337952
rect 271242 337940 271248 337952
rect 271242 337912 272150 337940
rect 271242 337900 271248 337912
rect 270374 337816 270402 337900
rect 270374 337776 270408 337816
rect 270402 337764 270408 337776
rect 270460 337764 270466 337816
rect 270092 337572 270218 337600
rect 270742 337612 270770 337900
rect 270908 337832 270914 337884
rect 270966 337832 270972 337884
rect 270742 337572 270776 337612
rect 270092 337560 270098 337572
rect 270770 337560 270776 337572
rect 270828 337560 270834 337612
rect 269178 337504 269212 337544
rect 269206 337492 269212 337504
rect 269264 337492 269270 337544
rect 270586 337492 270592 337544
rect 270644 337532 270650 337544
rect 270926 337532 270954 337832
rect 270644 337504 270954 337532
rect 270644 337492 270650 337504
rect 268160 337436 268838 337464
rect 268160 337424 268166 337436
rect 265860 337368 266124 337396
rect 271110 337396 271138 337900
rect 271552 337832 271558 337884
rect 271610 337832 271616 337884
rect 271828 337832 271834 337884
rect 271886 337832 271892 337884
rect 271230 337628 271236 337680
rect 271288 337668 271294 337680
rect 271570 337668 271598 337832
rect 271288 337640 271598 337668
rect 271288 337628 271294 337640
rect 271690 337628 271696 337680
rect 271748 337668 271754 337680
rect 271846 337668 271874 337832
rect 271748 337640 271874 337668
rect 271748 337628 271754 337640
rect 272122 337600 272150 337912
rect 272196 337900 272202 337952
rect 272254 337900 272260 337952
rect 272564 337900 272570 337952
rect 272622 337900 272628 337952
rect 272932 337900 272938 337952
rect 272990 337940 272996 337952
rect 272990 337900 273024 337940
rect 273116 337900 273122 337952
rect 273174 337900 273180 337952
rect 273760 337900 273766 337952
rect 273818 337900 273824 337952
rect 274128 337900 274134 337952
rect 274186 337900 274192 337952
rect 274220 337900 274226 337952
rect 274278 337900 274284 337952
rect 274312 337900 274318 337952
rect 274370 337900 274376 337952
rect 274496 337900 274502 337952
rect 274554 337900 274560 337952
rect 272214 337668 272242 337900
rect 272582 337680 272610 337900
rect 272996 337680 273024 337900
rect 272426 337668 272432 337680
rect 272214 337640 272432 337668
rect 272426 337628 272432 337640
rect 272484 337628 272490 337680
rect 272518 337628 272524 337680
rect 272576 337640 272610 337680
rect 272576 337628 272582 337640
rect 272978 337628 272984 337680
rect 273036 337628 273042 337680
rect 272334 337600 272340 337612
rect 272122 337572 272340 337600
rect 272334 337560 272340 337572
rect 272392 337560 272398 337612
rect 271966 337492 271972 337544
rect 272024 337532 272030 337544
rect 273134 337532 273162 337900
rect 273300 337832 273306 337884
rect 273358 337832 273364 337884
rect 273484 337832 273490 337884
rect 273542 337832 273548 337884
rect 273944 337872 273950 337884
rect 273732 337844 273950 337872
rect 272024 337504 273162 337532
rect 272024 337492 272030 337504
rect 273318 337464 273346 337832
rect 273502 337668 273530 337832
rect 273732 337816 273760 337844
rect 273944 337832 273950 337844
rect 274002 337832 274008 337884
rect 274036 337832 274042 337884
rect 274094 337832 274100 337884
rect 273714 337764 273720 337816
rect 273772 337764 273778 337816
rect 274054 337804 274082 337832
rect 274146 337816 274174 337900
rect 273916 337776 274082 337804
rect 273622 337668 273628 337680
rect 273502 337640 273628 337668
rect 273622 337628 273628 337640
rect 273680 337628 273686 337680
rect 273916 337532 273944 337776
rect 274128 337764 274134 337816
rect 274186 337764 274192 337816
rect 274238 337668 274266 337900
rect 274330 337816 274358 337900
rect 274514 337816 274542 337900
rect 274330 337776 274364 337816
rect 274358 337764 274364 337776
rect 274416 337764 274422 337816
rect 274450 337764 274456 337816
rect 274508 337776 274542 337816
rect 274606 337804 274634 337980
rect 274882 337980 275002 338008
rect 274606 337776 274680 337804
rect 274508 337764 274514 337776
rect 274542 337696 274548 337748
rect 274600 337736 274606 337748
rect 274652 337736 274680 337776
rect 274772 337764 274778 337816
rect 274830 337764 274836 337816
rect 274600 337708 274680 337736
rect 274600 337696 274606 337708
rect 274238 337640 274404 337668
rect 274082 337560 274088 337612
rect 274140 337600 274146 337612
rect 274266 337600 274272 337612
rect 274140 337572 274272 337600
rect 274140 337560 274146 337572
rect 274266 337560 274272 337572
rect 274324 337560 274330 337612
rect 273990 337532 273996 337544
rect 273916 337504 273996 337532
rect 273990 337492 273996 337504
rect 274048 337492 274054 337544
rect 274174 337492 274180 337544
rect 274232 337532 274238 337544
rect 274376 337532 274404 337640
rect 274232 337504 274404 337532
rect 274790 337532 274818 337764
rect 274882 337668 274910 337980
rect 274974 337952 275002 337980
rect 274956 337900 274962 337952
rect 275014 337900 275020 337952
rect 275508 337940 275514 337952
rect 275434 337912 275514 337940
rect 275048 337832 275054 337884
rect 275106 337832 275112 337884
rect 275140 337832 275146 337884
rect 275198 337872 275204 337884
rect 275198 337844 275370 337872
rect 275198 337832 275204 337844
rect 275066 337736 275094 337832
rect 275066 337708 275140 337736
rect 275002 337668 275008 337680
rect 274882 337640 275008 337668
rect 275002 337628 275008 337640
rect 275060 337628 275066 337680
rect 275112 337600 275140 337708
rect 275342 337612 275370 337844
rect 275434 337680 275462 337912
rect 275508 337900 275514 337912
rect 275566 337900 275572 337952
rect 275600 337872 275606 337884
rect 275572 337832 275606 337872
rect 275658 337832 275664 337884
rect 275572 337748 275600 337832
rect 275554 337696 275560 337748
rect 275612 337696 275618 337748
rect 275756 337680 275784 338184
rect 276354 337980 277118 338008
rect 276354 337952 276382 337980
rect 275876 337900 275882 337952
rect 275934 337900 275940 337952
rect 276152 337940 276158 337952
rect 276124 337900 276158 337940
rect 276210 337900 276216 337952
rect 276244 337900 276250 337952
rect 276302 337900 276308 337952
rect 276336 337900 276342 337952
rect 276394 337900 276400 337952
rect 276520 337900 276526 337952
rect 276578 337900 276584 337952
rect 276612 337900 276618 337952
rect 276670 337940 276676 337952
rect 276670 337900 276704 337940
rect 276796 337900 276802 337952
rect 276854 337900 276860 337952
rect 276888 337900 276894 337952
rect 276946 337900 276952 337952
rect 276980 337900 276986 337952
rect 277038 337900 277044 337952
rect 275434 337640 275468 337680
rect 275462 337628 275468 337640
rect 275520 337628 275526 337680
rect 275738 337628 275744 337680
rect 275796 337628 275802 337680
rect 275112 337572 275232 337600
rect 275342 337572 275376 337612
rect 274790 337504 275048 337532
rect 274232 337492 274238 337504
rect 274818 337464 274824 337476
rect 273318 337436 274824 337464
rect 274818 337424 274824 337436
rect 274876 337424 274882 337476
rect 274726 337396 274732 337408
rect 271110 337368 274732 337396
rect 265860 337356 265866 337368
rect 274726 337356 274732 337368
rect 274784 337356 274790 337408
rect 264204 337300 264376 337328
rect 264204 337288 264210 337300
rect 251634 337260 251640 337272
rect 244246 337232 251640 337260
rect 251634 337220 251640 337232
rect 251692 337220 251698 337272
rect 275020 337260 275048 337504
rect 275204 337340 275232 337572
rect 275370 337560 275376 337572
rect 275428 337560 275434 337612
rect 275894 337532 275922 337900
rect 275968 337832 275974 337884
rect 276026 337832 276032 337884
rect 275986 337612 276014 337832
rect 276124 337668 276152 337900
rect 276262 337816 276290 337900
rect 276198 337764 276204 337816
rect 276256 337776 276290 337816
rect 276256 337764 276262 337776
rect 276290 337668 276296 337680
rect 276124 337640 276296 337668
rect 276290 337628 276296 337640
rect 276348 337628 276354 337680
rect 275986 337572 276020 337612
rect 276014 337560 276020 337572
rect 276072 337560 276078 337612
rect 276538 337600 276566 337900
rect 276676 337680 276704 337900
rect 276814 337872 276842 337900
rect 276768 337844 276842 337872
rect 276658 337628 276664 337680
rect 276716 337628 276722 337680
rect 276538 337572 276704 337600
rect 276566 337532 276572 337544
rect 275894 337504 276572 337532
rect 276566 337492 276572 337504
rect 276624 337492 276630 337544
rect 276382 337424 276388 337476
rect 276440 337464 276446 337476
rect 276676 337464 276704 337572
rect 276440 337436 276704 337464
rect 276768 337464 276796 337844
rect 276906 337816 276934 337900
rect 276842 337764 276848 337816
rect 276900 337776 276934 337816
rect 276900 337764 276906 337776
rect 276998 337748 277026 337900
rect 276934 337696 276940 337748
rect 276992 337708 277026 337748
rect 276992 337696 276998 337708
rect 277090 337680 277118 337980
rect 277256 337900 277262 337952
rect 277314 337900 277320 337952
rect 277624 337900 277630 337952
rect 277682 337900 277688 337952
rect 277808 337900 277814 337952
rect 277866 337900 277872 337952
rect 277900 337900 277906 337952
rect 277958 337900 277964 337952
rect 277992 337900 277998 337952
rect 278050 337900 278056 337952
rect 278084 337900 278090 337952
rect 278142 337900 278148 337952
rect 278176 337900 278182 337952
rect 278234 337940 278240 337952
rect 278728 337940 278734 337952
rect 278234 337912 278636 337940
rect 278234 337900 278240 337912
rect 277026 337628 277032 337680
rect 277084 337640 277118 337680
rect 277084 337628 277090 337640
rect 277118 337492 277124 337544
rect 277176 337532 277182 337544
rect 277274 337532 277302 337900
rect 277642 337680 277670 337900
rect 277826 337872 277854 337900
rect 277780 337844 277854 337872
rect 277642 337640 277676 337680
rect 277670 337628 277676 337640
rect 277728 337628 277734 337680
rect 277780 337668 277808 337844
rect 277780 337640 277854 337668
rect 277176 337504 277302 337532
rect 277826 337544 277854 337640
rect 277918 337612 277946 337900
rect 278010 337816 278038 337900
rect 278102 337872 278130 337900
rect 278102 337844 278268 337872
rect 278010 337776 278044 337816
rect 278038 337764 278044 337776
rect 278096 337764 278102 337816
rect 277918 337572 277952 337612
rect 277946 337560 277952 337572
rect 278004 337560 278010 337612
rect 277826 337504 277860 337544
rect 277176 337492 277182 337504
rect 277854 337492 277860 337504
rect 277912 337492 277918 337544
rect 278240 337532 278268 337844
rect 278360 337804 278366 337816
rect 278332 337764 278366 337804
rect 278418 337764 278424 337816
rect 278332 337680 278360 337764
rect 278608 337680 278636 337912
rect 278700 337900 278734 337940
rect 278786 337900 278792 337952
rect 278912 337900 278918 337952
rect 278970 337900 278976 337952
rect 279004 337900 279010 337952
rect 279062 337900 279068 337952
rect 279096 337900 279102 337952
rect 279154 337900 279160 337952
rect 279188 337900 279194 337952
rect 279246 337900 279252 337952
rect 279280 337900 279286 337952
rect 279338 337940 279344 337952
rect 279464 337940 279470 337952
rect 279338 337900 279372 337940
rect 278700 337680 278728 337900
rect 278774 337764 278780 337816
rect 278832 337804 278838 337816
rect 278930 337804 278958 337900
rect 278832 337776 278958 337804
rect 278832 337764 278838 337776
rect 279022 337748 279050 337900
rect 278958 337696 278964 337748
rect 279016 337708 279050 337748
rect 279016 337696 279022 337708
rect 278314 337628 278320 337680
rect 278372 337628 278378 337680
rect 278590 337628 278596 337680
rect 278648 337628 278654 337680
rect 278682 337628 278688 337680
rect 278740 337628 278746 337680
rect 278866 337560 278872 337612
rect 278924 337600 278930 337612
rect 279114 337600 279142 337900
rect 278924 337572 279142 337600
rect 279206 337612 279234 337900
rect 279344 337612 279372 337900
rect 279436 337900 279470 337940
rect 279522 337900 279528 337952
rect 279556 337900 279562 337952
rect 279614 337900 279620 337952
rect 279648 337900 279654 337952
rect 279706 337900 279712 337952
rect 279832 337940 279838 337952
rect 279804 337900 279838 337940
rect 279890 337900 279896 337952
rect 280016 337900 280022 337952
rect 280074 337900 280080 337952
rect 279206 337572 279240 337612
rect 278924 337560 278930 337572
rect 279234 337560 279240 337572
rect 279292 337560 279298 337612
rect 279326 337560 279332 337612
rect 279384 337560 279390 337612
rect 279142 337532 279148 337544
rect 278240 337504 279148 337532
rect 279142 337492 279148 337504
rect 279200 337492 279206 337544
rect 278130 337464 278136 337476
rect 276768 337436 278136 337464
rect 276440 337424 276446 337436
rect 278130 337424 278136 337436
rect 278188 337424 278194 337476
rect 279436 337396 279464 337900
rect 279574 337872 279602 337900
rect 279528 337844 279602 337872
rect 279528 337748 279556 337844
rect 279666 337748 279694 337900
rect 279510 337696 279516 337748
rect 279568 337696 279574 337748
rect 279602 337696 279608 337748
rect 279660 337708 279694 337748
rect 279660 337696 279666 337708
rect 279804 337544 279832 337900
rect 280034 337872 280062 337900
rect 279896 337844 280062 337872
rect 279786 337492 279792 337544
rect 279844 337492 279850 337544
rect 279896 337476 279924 337844
rect 279970 337764 279976 337816
rect 280028 337804 280034 337816
rect 280126 337804 280154 338252
rect 430574 338240 430580 338252
rect 430632 338240 430638 338292
rect 448514 338212 448520 338224
rect 280218 338184 448520 338212
rect 280218 337952 280246 338184
rect 448514 338172 448520 338184
rect 448572 338172 448578 338224
rect 465074 338144 465080 338156
rect 281598 338116 465080 338144
rect 280200 337900 280206 337952
rect 280258 337900 280264 337952
rect 281028 337940 281034 337952
rect 280678 337912 281034 337940
rect 280476 337872 280482 337884
rect 280028 337776 280154 337804
rect 280356 337844 280482 337872
rect 280028 337764 280034 337776
rect 280356 337612 280384 337844
rect 280476 337832 280482 337844
rect 280534 337832 280540 337884
rect 280568 337832 280574 337884
rect 280626 337832 280632 337884
rect 280586 337680 280614 337832
rect 280522 337628 280528 337680
rect 280580 337640 280614 337680
rect 280580 337628 280586 337640
rect 280338 337560 280344 337612
rect 280396 337560 280402 337612
rect 280430 337560 280436 337612
rect 280488 337600 280494 337612
rect 280678 337600 280706 337912
rect 281028 337900 281034 337912
rect 281086 337900 281092 337952
rect 281396 337900 281402 337952
rect 281454 337900 281460 337952
rect 280936 337832 280942 337884
rect 280994 337832 281000 337884
rect 281120 337872 281126 337884
rect 281092 337832 281126 337872
rect 281178 337832 281184 337884
rect 281304 337832 281310 337884
rect 281362 337832 281368 337884
rect 280488 337572 280706 337600
rect 280954 337612 280982 337832
rect 281092 337748 281120 337832
rect 281212 337764 281218 337816
rect 281270 337764 281276 337816
rect 281074 337696 281080 337748
rect 281132 337696 281138 337748
rect 281230 337612 281258 337764
rect 280954 337572 280988 337612
rect 280488 337560 280494 337572
rect 280982 337560 280988 337572
rect 281040 337560 281046 337612
rect 281166 337560 281172 337612
rect 281224 337572 281258 337612
rect 281224 337560 281230 337572
rect 281322 337544 281350 337832
rect 281258 337492 281264 337544
rect 281316 337504 281350 337544
rect 281316 337492 281322 337504
rect 279878 337424 279884 337476
rect 279936 337424 279942 337476
rect 280798 337424 280804 337476
rect 280856 337464 280862 337476
rect 281414 337464 281442 337900
rect 281598 337884 281626 338116
rect 465074 338104 465080 338116
rect 465132 338104 465138 338156
rect 290918 338076 290924 338088
rect 287210 338048 290924 338076
rect 287210 337952 287238 338048
rect 290918 338036 290924 338048
rect 290976 338036 290982 338088
rect 290826 338008 290832 338020
rect 289878 337980 290832 338008
rect 281764 337900 281770 337952
rect 281822 337900 281828 337952
rect 282132 337900 282138 337952
rect 282190 337900 282196 337952
rect 282224 337900 282230 337952
rect 282282 337900 282288 337952
rect 282960 337900 282966 337952
rect 283018 337900 283024 337952
rect 283972 337900 283978 337952
rect 284030 337900 284036 337952
rect 284340 337900 284346 337952
rect 284398 337900 284404 337952
rect 284524 337900 284530 337952
rect 284582 337900 284588 337952
rect 285260 337940 285266 337952
rect 284864 337912 285266 337940
rect 281580 337832 281586 337884
rect 281638 337832 281644 337884
rect 281782 337736 281810 337900
rect 281948 337832 281954 337884
rect 282006 337832 282012 337884
rect 281552 337708 281810 337736
rect 281552 337680 281580 337708
rect 281534 337628 281540 337680
rect 281592 337628 281598 337680
rect 281626 337560 281632 337612
rect 281684 337600 281690 337612
rect 281966 337600 281994 337832
rect 282150 337748 282178 337900
rect 282086 337696 282092 337748
rect 282144 337708 282178 337748
rect 282144 337696 282150 337708
rect 282242 337680 282270 337900
rect 282592 337832 282598 337884
rect 282650 337832 282656 337884
rect 282868 337832 282874 337884
rect 282926 337832 282932 337884
rect 282242 337640 282276 337680
rect 282270 337628 282276 337640
rect 282328 337628 282334 337680
rect 281684 337572 281994 337600
rect 282610 337612 282638 337832
rect 282610 337572 282644 337612
rect 281684 337560 281690 337572
rect 282638 337560 282644 337572
rect 282696 337560 282702 337612
rect 280856 337436 281442 337464
rect 280856 337424 280862 337436
rect 280062 337396 280068 337408
rect 279436 337368 280068 337396
rect 280062 337356 280068 337368
rect 280120 337356 280126 337408
rect 281442 337356 281448 337408
rect 281500 337356 281506 337408
rect 275186 337288 275192 337340
rect 275244 337288 275250 337340
rect 281460 337328 281488 337356
rect 282454 337328 282460 337340
rect 281460 337300 282460 337328
rect 282454 337288 282460 337300
rect 282512 337288 282518 337340
rect 275094 337260 275100 337272
rect 275020 337232 275100 337260
rect 275094 337220 275100 337232
rect 275152 337220 275158 337272
rect 280246 337220 280252 337272
rect 280304 337260 280310 337272
rect 281442 337260 281448 337272
rect 280304 337232 281448 337260
rect 280304 337220 280310 337232
rect 281442 337220 281448 337232
rect 281500 337220 281506 337272
rect 281902 337220 281908 337272
rect 281960 337260 281966 337272
rect 282886 337260 282914 337832
rect 281960 337232 282914 337260
rect 282978 337260 283006 337900
rect 283328 337832 283334 337884
rect 283386 337832 283392 337884
rect 283604 337832 283610 337884
rect 283662 337832 283668 337884
rect 283144 337804 283150 337816
rect 283116 337764 283150 337804
rect 283202 337764 283208 337816
rect 283116 337680 283144 337764
rect 283098 337628 283104 337680
rect 283156 337628 283162 337680
rect 283346 337544 283374 337832
rect 283622 337600 283650 337832
rect 283990 337816 284018 337900
rect 283926 337764 283932 337816
rect 283984 337776 284018 337816
rect 283984 337764 283990 337776
rect 284064 337764 284070 337816
rect 284122 337764 284128 337816
rect 284248 337764 284254 337816
rect 284306 337764 284312 337816
rect 284082 337680 284110 337764
rect 284018 337628 284024 337680
rect 284076 337640 284110 337680
rect 284076 337628 284082 337640
rect 283484 337572 283650 337600
rect 283484 337544 283512 337572
rect 284266 337544 284294 337764
rect 284358 337612 284386 337900
rect 284542 337748 284570 337900
rect 284616 337832 284622 337884
rect 284674 337832 284680 337884
rect 284708 337832 284714 337884
rect 284766 337832 284772 337884
rect 284478 337696 284484 337748
rect 284536 337708 284570 337748
rect 284536 337696 284542 337708
rect 284634 337680 284662 337832
rect 284570 337628 284576 337680
rect 284628 337640 284662 337680
rect 284628 337628 284634 337640
rect 284726 337612 284754 337832
rect 284358 337572 284392 337612
rect 284386 337560 284392 337572
rect 284444 337560 284450 337612
rect 284662 337560 284668 337612
rect 284720 337572 284754 337612
rect 284720 337560 284726 337572
rect 283282 337492 283288 337544
rect 283340 337504 283374 337544
rect 283340 337492 283346 337504
rect 283466 337492 283472 337544
rect 283524 337492 283530 337544
rect 284202 337492 284208 337544
rect 284260 337504 284294 337544
rect 284260 337492 284266 337504
rect 284864 337464 284892 337912
rect 285260 337900 285266 337912
rect 285318 337900 285324 337952
rect 286456 337900 286462 337952
rect 286514 337900 286520 337952
rect 286548 337900 286554 337952
rect 286606 337900 286612 337952
rect 286640 337900 286646 337952
rect 286698 337940 286704 337952
rect 286698 337900 286732 337940
rect 287008 337900 287014 337952
rect 287066 337900 287072 337952
rect 287192 337900 287198 337952
rect 287250 337900 287256 337952
rect 287376 337900 287382 337952
rect 287434 337900 287440 337952
rect 287560 337900 287566 337952
rect 287618 337900 287624 337952
rect 287652 337900 287658 337952
rect 287710 337900 287716 337952
rect 287928 337900 287934 337952
rect 287986 337900 287992 337952
rect 288020 337900 288026 337952
rect 288078 337900 288084 337952
rect 288204 337900 288210 337952
rect 288262 337900 288268 337952
rect 288572 337900 288578 337952
rect 288630 337900 288636 337952
rect 289216 337940 289222 337952
rect 289188 337900 289222 337940
rect 289274 337900 289280 337952
rect 289676 337900 289682 337952
rect 289734 337900 289740 337952
rect 285168 337832 285174 337884
rect 285226 337832 285232 337884
rect 285352 337832 285358 337884
rect 285410 337832 285416 337884
rect 285444 337832 285450 337884
rect 285502 337832 285508 337884
rect 285536 337832 285542 337884
rect 285594 337832 285600 337884
rect 286088 337832 286094 337884
rect 286146 337832 286152 337884
rect 285186 337544 285214 337832
rect 285370 337736 285398 337832
rect 285324 337708 285398 337736
rect 285324 337680 285352 337708
rect 285462 337680 285490 337832
rect 285306 337628 285312 337680
rect 285364 337628 285370 337680
rect 285398 337628 285404 337680
rect 285456 337640 285490 337680
rect 285456 337628 285462 337640
rect 285122 337492 285128 337544
rect 285180 337504 285214 337544
rect 285180 337492 285186 337504
rect 285030 337464 285036 337476
rect 284864 337436 285036 337464
rect 285030 337424 285036 337436
rect 285088 337424 285094 337476
rect 285214 337424 285220 337476
rect 285272 337464 285278 337476
rect 285554 337464 285582 337832
rect 286106 337600 286134 337832
rect 286474 337816 286502 337900
rect 286566 337872 286594 337900
rect 286566 337844 286640 337872
rect 286612 337816 286640 337844
rect 286474 337776 286508 337816
rect 286502 337764 286508 337776
rect 286560 337764 286566 337816
rect 286594 337764 286600 337816
rect 286652 337764 286658 337816
rect 286704 337680 286732 337900
rect 286824 337764 286830 337816
rect 286882 337764 286888 337816
rect 287026 337804 287054 337900
rect 287238 337804 287244 337816
rect 287026 337776 287244 337804
rect 287238 337764 287244 337776
rect 287296 337764 287302 337816
rect 286842 337680 286870 337764
rect 286686 337628 286692 337680
rect 286744 337628 286750 337680
rect 286842 337640 286876 337680
rect 286870 337628 286876 337640
rect 286928 337628 286934 337680
rect 286226 337600 286232 337612
rect 286106 337572 286232 337600
rect 286226 337560 286232 337572
rect 286284 337560 286290 337612
rect 287394 337600 287422 337900
rect 287578 337816 287606 337900
rect 287514 337764 287520 337816
rect 287572 337776 287606 337816
rect 287572 337764 287578 337776
rect 287670 337680 287698 337900
rect 287836 337764 287842 337816
rect 287894 337764 287900 337816
rect 287854 337680 287882 337764
rect 287606 337628 287612 337680
rect 287664 337640 287698 337680
rect 287664 337628 287670 337640
rect 287790 337628 287796 337680
rect 287848 337640 287882 337680
rect 287848 337628 287854 337640
rect 287698 337600 287704 337612
rect 287394 337572 287704 337600
rect 287698 337560 287704 337572
rect 287756 337560 287762 337612
rect 287146 337492 287152 337544
rect 287204 337532 287210 337544
rect 287606 337532 287612 337544
rect 287204 337504 287612 337532
rect 287204 337492 287210 337504
rect 287606 337492 287612 337504
rect 287664 337492 287670 337544
rect 285272 337436 285582 337464
rect 285272 337424 285278 337436
rect 286962 337424 286968 337476
rect 287020 337464 287026 337476
rect 287946 337464 287974 337900
rect 288038 337612 288066 337900
rect 288222 337816 288250 337900
rect 288296 337832 288302 337884
rect 288354 337832 288360 337884
rect 288204 337764 288210 337816
rect 288262 337764 288268 337816
rect 288314 337680 288342 337832
rect 288590 337804 288618 337900
rect 288664 337832 288670 337884
rect 288722 337872 288728 337884
rect 288722 337844 289124 337872
rect 288722 337832 288728 337844
rect 288848 337804 288854 337816
rect 288590 337776 288664 337804
rect 288636 337748 288664 337776
rect 288820 337764 288854 337804
rect 288906 337764 288912 337816
rect 288618 337696 288624 337748
rect 288676 337696 288682 337748
rect 288250 337628 288256 337680
rect 288308 337640 288342 337680
rect 288308 337628 288314 337640
rect 288038 337572 288072 337612
rect 288066 337560 288072 337572
rect 288124 337560 288130 337612
rect 288820 337544 288848 337764
rect 288940 337696 288946 337748
rect 288998 337696 289004 337748
rect 288802 337492 288808 337544
rect 288860 337492 288866 337544
rect 287020 337436 287974 337464
rect 287020 337424 287026 337436
rect 288434 337424 288440 337476
rect 288492 337464 288498 337476
rect 288958 337464 288986 337696
rect 289096 337612 289124 337844
rect 289188 337680 289216 337900
rect 289308 337764 289314 337816
rect 289366 337764 289372 337816
rect 289400 337764 289406 337816
rect 289458 337764 289464 337816
rect 289694 337804 289722 337900
rect 289878 337884 289906 337980
rect 290826 337968 290832 337980
rect 290884 337968 290890 338020
rect 290044 337900 290050 337952
rect 290102 337900 290108 337952
rect 290228 337900 290234 337952
rect 290286 337900 290292 337952
rect 290320 337900 290326 337952
rect 290378 337940 290384 337952
rect 290378 337900 290412 337940
rect 290504 337900 290510 337952
rect 290562 337900 290568 337952
rect 289860 337832 289866 337884
rect 289918 337832 289924 337884
rect 289952 337832 289958 337884
rect 290010 337832 290016 337884
rect 289694 337776 289768 337804
rect 289170 337628 289176 337680
rect 289228 337628 289234 337680
rect 289326 337612 289354 337764
rect 289418 337736 289446 337764
rect 289630 337736 289636 337748
rect 289418 337708 289636 337736
rect 289630 337696 289636 337708
rect 289688 337696 289694 337748
rect 289740 337680 289768 337776
rect 289970 337680 289998 337832
rect 290062 337748 290090 337900
rect 290246 337872 290274 337900
rect 290246 337844 290320 337872
rect 290062 337708 290096 337748
rect 290090 337696 290096 337708
rect 290148 337696 290154 337748
rect 289722 337628 289728 337680
rect 289780 337628 289786 337680
rect 289906 337628 289912 337680
rect 289964 337640 289998 337680
rect 290292 337668 290320 337844
rect 290384 337680 290412 337900
rect 290522 337680 290550 337900
rect 290062 337640 290320 337668
rect 289964 337628 289970 337640
rect 289078 337560 289084 337612
rect 289136 337560 289142 337612
rect 289326 337572 289360 337612
rect 289354 337560 289360 337572
rect 289412 337560 289418 337612
rect 289814 337560 289820 337612
rect 289872 337600 289878 337612
rect 290062 337600 290090 337640
rect 290366 337628 290372 337680
rect 290424 337628 290430 337680
rect 290458 337628 290464 337680
rect 290516 337640 290550 337680
rect 290516 337628 290522 337640
rect 289872 337572 290090 337600
rect 289872 337560 289878 337572
rect 288492 337436 288986 337464
rect 288492 337424 288498 337436
rect 283742 337396 283748 337408
rect 283576 337368 283748 337396
rect 283576 337340 283604 337368
rect 283742 337356 283748 337368
rect 283800 337356 283806 337408
rect 287606 337356 287612 337408
rect 287664 337396 287670 337408
rect 346578 337396 346584 337408
rect 287664 337368 346584 337396
rect 287664 337356 287670 337368
rect 346578 337356 346584 337368
rect 346636 337356 346642 337408
rect 283558 337288 283564 337340
rect 283616 337288 283622 337340
rect 288066 337288 288072 337340
rect 288124 337328 288130 337340
rect 346670 337328 346676 337340
rect 288124 337300 346676 337328
rect 288124 337288 288130 337300
rect 346670 337288 346676 337300
rect 346728 337288 346734 337340
rect 283742 337260 283748 337272
rect 282978 337232 283748 337260
rect 281960 337220 281966 337232
rect 283742 337220 283748 337232
rect 283800 337220 283806 337272
rect 285582 337220 285588 337272
rect 285640 337260 285646 337272
rect 345658 337260 345664 337272
rect 285640 337232 345664 337260
rect 285640 337220 285646 337232
rect 345658 337220 345664 337232
rect 345716 337220 345722 337272
rect 227714 337152 227720 337204
rect 227772 337192 227778 337204
rect 263134 337192 263140 337204
rect 227772 337164 263140 337192
rect 227772 337152 227778 337164
rect 263134 337152 263140 337164
rect 263192 337152 263198 337204
rect 271874 337152 271880 337204
rect 271932 337192 271938 337204
rect 346486 337192 346492 337204
rect 271932 337164 273254 337192
rect 271932 337152 271938 337164
rect 218054 337084 218060 337136
rect 218112 337124 218118 337136
rect 262214 337124 262220 337136
rect 218112 337096 262220 337124
rect 218112 337084 218118 337096
rect 262214 337084 262220 337096
rect 262272 337084 262278 337136
rect 273226 337124 273254 337164
rect 274836 337164 346492 337192
rect 274836 337124 274864 337164
rect 346486 337152 346492 337164
rect 346544 337152 346550 337204
rect 273226 337096 274864 337124
rect 275738 337084 275744 337136
rect 275796 337124 275802 337136
rect 343910 337124 343916 337136
rect 275796 337096 343916 337124
rect 275796 337084 275802 337096
rect 343910 337084 343916 337096
rect 343968 337084 343974 337136
rect 165614 337016 165620 337068
rect 165672 337056 165678 337068
rect 248966 337056 248972 337068
rect 165672 337028 248972 337056
rect 165672 337016 165678 337028
rect 248966 337016 248972 337028
rect 249024 337016 249030 337068
rect 250162 337016 250168 337068
rect 250220 337056 250226 337068
rect 250622 337056 250628 337068
rect 250220 337028 250628 337056
rect 250220 337016 250226 337028
rect 250622 337016 250628 337028
rect 250680 337016 250686 337068
rect 346394 337056 346400 337068
rect 276032 337028 346400 337056
rect 161474 336948 161480 337000
rect 161532 336988 161538 337000
rect 257890 336988 257896 337000
rect 161532 336960 257896 336988
rect 161532 336948 161538 336960
rect 257890 336948 257896 336960
rect 257948 336948 257954 337000
rect 270034 336948 270040 337000
rect 270092 336988 270098 337000
rect 276032 336988 276060 337028
rect 346394 337016 346400 337028
rect 346452 337016 346458 337068
rect 270092 336960 276060 336988
rect 270092 336948 270098 336960
rect 276106 336948 276112 337000
rect 276164 336988 276170 337000
rect 394694 336988 394700 337000
rect 276164 336960 394700 336988
rect 276164 336948 276170 336960
rect 394694 336948 394700 336960
rect 394752 336948 394758 337000
rect 241422 336880 241428 336932
rect 241480 336920 241486 336932
rect 249794 336920 249800 336932
rect 241480 336892 249800 336920
rect 241480 336880 241486 336892
rect 249794 336880 249800 336892
rect 249852 336880 249858 336932
rect 267274 336920 267280 336932
rect 253906 336892 267280 336920
rect 240042 336812 240048 336864
rect 240100 336852 240106 336864
rect 253906 336852 253934 336892
rect 267274 336880 267280 336892
rect 267332 336880 267338 336932
rect 272426 336880 272432 336932
rect 272484 336920 272490 336932
rect 272484 336892 274634 336920
rect 272484 336880 272490 336892
rect 240100 336824 253934 336852
rect 240100 336812 240106 336824
rect 273622 336812 273628 336864
rect 273680 336812 273686 336864
rect 234614 336744 234620 336796
rect 234672 336784 234678 336796
rect 263686 336784 263692 336796
rect 234672 336756 263692 336784
rect 234672 336744 234678 336756
rect 263686 336744 263692 336756
rect 263744 336744 263750 336796
rect 273640 336784 273668 336812
rect 273640 336756 273760 336784
rect 242342 336676 242348 336728
rect 242400 336716 242406 336728
rect 246758 336716 246764 336728
rect 242400 336688 246764 336716
rect 242400 336676 242406 336688
rect 246758 336676 246764 336688
rect 246816 336676 246822 336728
rect 256418 336676 256424 336728
rect 256476 336716 256482 336728
rect 268194 336716 268200 336728
rect 256476 336688 268200 336716
rect 256476 336676 256482 336688
rect 268194 336676 268200 336688
rect 268252 336676 268258 336728
rect 244182 336608 244188 336660
rect 244240 336648 244246 336660
rect 244240 336608 244274 336648
rect 248414 336608 248420 336660
rect 248472 336648 248478 336660
rect 260926 336648 260932 336660
rect 248472 336620 260932 336648
rect 248472 336608 248478 336620
rect 260926 336608 260932 336620
rect 260984 336608 260990 336660
rect 273732 336648 273760 336756
rect 274606 336716 274634 336892
rect 277210 336880 277216 336932
rect 277268 336920 277274 336932
rect 408494 336920 408500 336932
rect 277268 336892 408500 336920
rect 277268 336880 277274 336892
rect 408494 336880 408500 336892
rect 408552 336880 408558 336932
rect 280338 336812 280344 336864
rect 280396 336852 280402 336864
rect 451274 336852 451280 336864
rect 280396 336824 451280 336852
rect 280396 336812 280402 336824
rect 451274 336812 451280 336824
rect 451332 336812 451338 336864
rect 280246 336744 280252 336796
rect 280304 336784 280310 336796
rect 281166 336784 281172 336796
rect 280304 336756 281172 336784
rect 280304 336744 280310 336756
rect 281166 336744 281172 336756
rect 281224 336744 281230 336796
rect 281718 336744 281724 336796
rect 281776 336784 281782 336796
rect 282546 336784 282552 336796
rect 281776 336756 282552 336784
rect 281776 336744 281782 336756
rect 282546 336744 282552 336756
rect 282604 336744 282610 336796
rect 292850 336744 292856 336796
rect 292908 336784 292914 336796
rect 557534 336784 557540 336796
rect 292908 336756 557540 336784
rect 292908 336744 292914 336756
rect 557534 336744 557540 336756
rect 557592 336744 557598 336796
rect 285582 336716 285588 336728
rect 274606 336688 285588 336716
rect 285582 336676 285588 336688
rect 285640 336676 285646 336728
rect 287238 336676 287244 336728
rect 287296 336716 287302 336728
rect 291194 336716 291200 336728
rect 287296 336688 291200 336716
rect 287296 336676 287302 336688
rect 291194 336676 291200 336688
rect 291252 336676 291258 336728
rect 277302 336648 277308 336660
rect 273732 336620 277308 336648
rect 277302 336608 277308 336620
rect 277360 336608 277366 336660
rect 287606 336648 287612 336660
rect 277412 336620 287612 336648
rect 244246 336580 244274 336608
rect 264974 336580 264980 336592
rect 244246 336552 264980 336580
rect 264974 336540 264980 336552
rect 265032 336540 265038 336592
rect 274726 336540 274732 336592
rect 274784 336580 274790 336592
rect 277412 336580 277440 336620
rect 287606 336608 287612 336620
rect 287664 336608 287670 336660
rect 274784 336552 277440 336580
rect 274784 336540 274790 336552
rect 279786 336540 279792 336592
rect 279844 336580 279850 336592
rect 285306 336580 285312 336592
rect 279844 336552 285312 336580
rect 279844 336540 279850 336552
rect 285306 336540 285312 336552
rect 285364 336540 285370 336592
rect 287238 336540 287244 336592
rect 287296 336580 287302 336592
rect 293402 336580 293408 336592
rect 287296 336552 293408 336580
rect 287296 336540 287302 336552
rect 293402 336540 293408 336552
rect 293460 336540 293466 336592
rect 224954 336472 224960 336524
rect 225012 336512 225018 336524
rect 262306 336512 262312 336524
rect 225012 336484 262312 336512
rect 225012 336472 225018 336484
rect 262306 336472 262312 336484
rect 262364 336472 262370 336524
rect 278682 336472 278688 336524
rect 278740 336512 278746 336524
rect 287882 336512 287888 336524
rect 278740 336484 287888 336512
rect 278740 336472 278746 336484
rect 287882 336472 287888 336484
rect 287940 336472 287946 336524
rect 196618 336404 196624 336456
rect 196676 336444 196682 336456
rect 247770 336444 247776 336456
rect 196676 336416 247776 336444
rect 196676 336404 196682 336416
rect 247770 336404 247776 336416
rect 247828 336404 247834 336456
rect 277394 336404 277400 336456
rect 277452 336444 277458 336456
rect 293218 336444 293224 336456
rect 277452 336416 293224 336444
rect 277452 336404 277458 336416
rect 293218 336404 293224 336416
rect 293276 336404 293282 336456
rect 200758 336336 200764 336388
rect 200816 336376 200822 336388
rect 248598 336376 248604 336388
rect 200816 336348 248604 336376
rect 200816 336336 200822 336348
rect 248598 336336 248604 336348
rect 248656 336336 248662 336388
rect 249794 336336 249800 336388
rect 249852 336376 249858 336388
rect 249852 336348 263594 336376
rect 249852 336336 249858 336348
rect 188338 336268 188344 336320
rect 188396 336308 188402 336320
rect 247494 336308 247500 336320
rect 188396 336280 247500 336308
rect 188396 336268 188402 336280
rect 247494 336268 247500 336280
rect 247552 336268 247558 336320
rect 255498 336268 255504 336320
rect 255556 336308 255562 336320
rect 256602 336308 256608 336320
rect 255556 336280 256608 336308
rect 255556 336268 255562 336280
rect 256602 336268 256608 336280
rect 256660 336268 256666 336320
rect 258442 336268 258448 336320
rect 258500 336308 258506 336320
rect 259178 336308 259184 336320
rect 258500 336280 259184 336308
rect 258500 336268 258506 336280
rect 259178 336268 259184 336280
rect 259236 336268 259242 336320
rect 259730 336268 259736 336320
rect 259788 336308 259794 336320
rect 260282 336308 260288 336320
rect 259788 336280 260288 336308
rect 259788 336268 259794 336280
rect 260282 336268 260288 336280
rect 260340 336268 260346 336320
rect 182174 336200 182180 336252
rect 182232 336240 182238 336252
rect 248966 336240 248972 336252
rect 182232 336212 248972 336240
rect 182232 336200 182238 336212
rect 248966 336200 248972 336212
rect 249024 336200 249030 336252
rect 253566 336200 253572 336252
rect 253624 336240 253630 336252
rect 262674 336240 262680 336252
rect 253624 336212 262680 336240
rect 253624 336200 253630 336212
rect 262674 336200 262680 336212
rect 262732 336200 262738 336252
rect 263566 336240 263594 336348
rect 276014 336336 276020 336388
rect 276072 336376 276078 336388
rect 291930 336376 291936 336388
rect 276072 336348 291936 336376
rect 276072 336336 276078 336348
rect 291930 336336 291936 336348
rect 291988 336336 291994 336388
rect 280706 336268 280712 336320
rect 280764 336308 280770 336320
rect 346762 336308 346768 336320
rect 280764 336280 346768 336308
rect 280764 336268 280770 336280
rect 346762 336268 346768 336280
rect 346820 336268 346826 336320
rect 266262 336240 266268 336252
rect 263566 336212 266268 336240
rect 266262 336200 266268 336212
rect 266320 336200 266326 336252
rect 270402 336200 270408 336252
rect 270460 336240 270466 336252
rect 279878 336240 279884 336252
rect 270460 336212 279884 336240
rect 270460 336200 270466 336212
rect 279878 336200 279884 336212
rect 279936 336200 279942 336252
rect 281534 336200 281540 336252
rect 281592 336240 281598 336252
rect 467834 336240 467840 336252
rect 281592 336212 467840 336240
rect 281592 336200 281598 336212
rect 467834 336200 467840 336212
rect 467892 336200 467898 336252
rect 160094 336132 160100 336184
rect 160152 336172 160158 336184
rect 257798 336172 257804 336184
rect 160152 336144 257804 336172
rect 160152 336132 160158 336144
rect 257798 336132 257804 336144
rect 257856 336132 257862 336184
rect 257890 336132 257896 336184
rect 257948 336172 257954 336184
rect 264238 336172 264244 336184
rect 257948 336144 264244 336172
rect 257948 336132 257954 336144
rect 264238 336132 264244 336144
rect 264296 336132 264302 336184
rect 277578 336132 277584 336184
rect 277636 336172 277642 336184
rect 278958 336172 278964 336184
rect 277636 336144 278964 336172
rect 277636 336132 277642 336144
rect 278958 336132 278964 336144
rect 279016 336132 279022 336184
rect 281350 336132 281356 336184
rect 281408 336172 281414 336184
rect 283190 336172 283196 336184
rect 281408 336144 283196 336172
rect 281408 336132 281414 336144
rect 283190 336132 283196 336144
rect 283248 336132 283254 336184
rect 283742 336132 283748 336184
rect 283800 336172 283806 336184
rect 483014 336172 483020 336184
rect 283800 336144 483020 336172
rect 283800 336132 283806 336144
rect 483014 336132 483020 336144
rect 483072 336132 483078 336184
rect 128354 336064 128360 336116
rect 128412 336104 128418 336116
rect 255314 336104 255320 336116
rect 128412 336076 255320 336104
rect 128412 336064 128418 336076
rect 255314 336064 255320 336076
rect 255372 336064 255378 336116
rect 267734 336104 267740 336116
rect 255424 336076 267740 336104
rect 125594 335996 125600 336048
rect 125652 336036 125658 336048
rect 255038 336036 255044 336048
rect 125652 336008 255044 336036
rect 125652 335996 125658 336008
rect 255038 335996 255044 336008
rect 255096 335996 255102 336048
rect 242434 335928 242440 335980
rect 242492 335968 242498 335980
rect 253290 335968 253296 335980
rect 242492 335940 253296 335968
rect 242492 335928 242498 335940
rect 253290 335928 253296 335940
rect 253348 335928 253354 335980
rect 255314 335928 255320 335980
rect 255372 335968 255378 335980
rect 255424 335968 255452 336076
rect 267734 336064 267740 336076
rect 267792 336064 267798 336116
rect 281534 336064 281540 336116
rect 281592 336104 281598 336116
rect 282270 336104 282276 336116
rect 281592 336076 282276 336104
rect 281592 336064 281598 336076
rect 282270 336064 282276 336076
rect 282328 336064 282334 336116
rect 284386 336064 284392 336116
rect 284444 336104 284450 336116
rect 500954 336104 500960 336116
rect 284444 336076 500960 336104
rect 284444 336064 284450 336076
rect 500954 336064 500960 336076
rect 501012 336064 501018 336116
rect 256418 335996 256424 336048
rect 256476 336036 256482 336048
rect 273254 336036 273260 336048
rect 256476 336008 273260 336036
rect 256476 335996 256482 336008
rect 273254 335996 273260 336008
rect 273312 335996 273318 336048
rect 287054 335996 287060 336048
rect 287112 336036 287118 336048
rect 536834 336036 536840 336048
rect 287112 336008 536840 336036
rect 287112 335996 287118 336008
rect 536834 335996 536840 336008
rect 536892 335996 536898 336048
rect 255372 335940 255452 335968
rect 255372 335928 255378 335940
rect 259178 335928 259184 335980
rect 259236 335968 259242 335980
rect 268470 335968 268476 335980
rect 259236 335940 268476 335968
rect 259236 335928 259242 335940
rect 268470 335928 268476 335940
rect 268528 335928 268534 335980
rect 269942 335928 269948 335980
rect 270000 335968 270006 335980
rect 270218 335968 270224 335980
rect 270000 335940 270224 335968
rect 270000 335928 270006 335940
rect 270218 335928 270224 335940
rect 270276 335928 270282 335980
rect 278130 335928 278136 335980
rect 278188 335968 278194 335980
rect 292114 335968 292120 335980
rect 278188 335940 292120 335968
rect 278188 335928 278194 335940
rect 292114 335928 292120 335940
rect 292172 335928 292178 335980
rect 243722 335860 243728 335912
rect 243780 335900 243786 335912
rect 251910 335900 251916 335912
rect 243780 335872 251916 335900
rect 243780 335860 243786 335872
rect 251910 335860 251916 335872
rect 251968 335860 251974 335912
rect 260006 335860 260012 335912
rect 260064 335900 260070 335912
rect 260282 335900 260288 335912
rect 260064 335872 260288 335900
rect 260064 335860 260070 335872
rect 260282 335860 260288 335872
rect 260340 335860 260346 335912
rect 262674 335860 262680 335912
rect 262732 335900 262738 335912
rect 262950 335900 262956 335912
rect 262732 335872 262956 335900
rect 262732 335860 262738 335872
rect 262950 335860 262956 335872
rect 263008 335860 263014 335912
rect 277394 335860 277400 335912
rect 277452 335900 277458 335912
rect 277762 335900 277768 335912
rect 277452 335872 277768 335900
rect 277452 335860 277458 335872
rect 277762 335860 277768 335872
rect 277820 335860 277826 335912
rect 278590 335860 278596 335912
rect 278648 335900 278654 335912
rect 287238 335900 287244 335912
rect 278648 335872 287244 335900
rect 278648 335860 278654 335872
rect 287238 335860 287244 335872
rect 287296 335860 287302 335912
rect 287882 335860 287888 335912
rect 287940 335900 287946 335912
rect 293310 335900 293316 335912
rect 287940 335872 293316 335900
rect 287940 335860 287946 335872
rect 293310 335860 293316 335872
rect 293368 335860 293374 335912
rect 242158 335792 242164 335844
rect 242216 335832 242222 335844
rect 248414 335832 248420 335844
rect 242216 335804 248420 335832
rect 242216 335792 242222 335804
rect 248414 335792 248420 335804
rect 248472 335792 248478 335844
rect 248966 335792 248972 335844
rect 249024 335832 249030 335844
rect 259454 335832 259460 335844
rect 249024 335804 259460 335832
rect 249024 335792 249030 335804
rect 259454 335792 259460 335804
rect 259512 335792 259518 335844
rect 279326 335792 279332 335844
rect 279384 335832 279390 335844
rect 293494 335832 293500 335844
rect 279384 335804 293500 335832
rect 279384 335792 279390 335804
rect 293494 335792 293500 335804
rect 293552 335792 293558 335844
rect 243906 335724 243912 335776
rect 243964 335764 243970 335776
rect 252462 335764 252468 335776
rect 243964 335736 252468 335764
rect 243964 335724 243970 335736
rect 252462 335724 252468 335736
rect 252520 335724 252526 335776
rect 255774 335724 255780 335776
rect 255832 335764 255838 335776
rect 255958 335764 255964 335776
rect 255832 335736 255964 335764
rect 255832 335724 255838 335736
rect 255958 335724 255964 335736
rect 256016 335724 256022 335776
rect 261294 335724 261300 335776
rect 261352 335764 261358 335776
rect 261570 335764 261576 335776
rect 261352 335736 261576 335764
rect 261352 335724 261358 335736
rect 261570 335724 261576 335736
rect 261628 335724 261634 335776
rect 283190 335724 283196 335776
rect 283248 335764 283254 335776
rect 294598 335764 294604 335776
rect 283248 335736 294604 335764
rect 283248 335724 283254 335736
rect 294598 335724 294604 335736
rect 294656 335724 294662 335776
rect 248966 335656 248972 335708
rect 249024 335696 249030 335708
rect 261754 335696 261760 335708
rect 249024 335668 261760 335696
rect 249024 335656 249030 335668
rect 261754 335656 261760 335668
rect 261812 335656 261818 335708
rect 273162 335656 273168 335708
rect 273220 335696 273226 335708
rect 288066 335696 288072 335708
rect 273220 335668 288072 335696
rect 273220 335656 273226 335668
rect 288066 335656 288072 335668
rect 288124 335656 288130 335708
rect 251910 335588 251916 335640
rect 251968 335628 251974 335640
rect 255866 335628 255872 335640
rect 251968 335600 255872 335628
rect 251968 335588 251974 335600
rect 255866 335588 255872 335600
rect 255924 335588 255930 335640
rect 277302 335588 277308 335640
rect 277360 335628 277366 335640
rect 281350 335628 281356 335640
rect 277360 335600 281356 335628
rect 277360 335588 277366 335600
rect 281350 335588 281356 335600
rect 281408 335588 281414 335640
rect 292022 335628 292028 335640
rect 285646 335600 292028 335628
rect 252462 335520 252468 335572
rect 252520 335560 252526 335572
rect 252520 335532 253934 335560
rect 252520 335520 252526 335532
rect 253906 335492 253934 335532
rect 261570 335520 261576 335572
rect 261628 335560 261634 335572
rect 265342 335560 265348 335572
rect 261628 335532 265348 335560
rect 261628 335520 261634 335532
rect 265342 335520 265348 335532
rect 265400 335520 265406 335572
rect 276198 335520 276204 335572
rect 276256 335560 276262 335572
rect 285646 335560 285674 335600
rect 292022 335588 292028 335600
rect 292080 335588 292086 335640
rect 276256 335532 285674 335560
rect 276256 335520 276262 335532
rect 258166 335492 258172 335504
rect 253906 335464 258172 335492
rect 258166 335452 258172 335464
rect 258224 335452 258230 335504
rect 274910 335452 274916 335504
rect 274968 335492 274974 335504
rect 281810 335492 281816 335504
rect 274968 335464 281816 335492
rect 274968 335452 274974 335464
rect 281810 335452 281816 335464
rect 281868 335452 281874 335504
rect 252186 335384 252192 335436
rect 252244 335424 252250 335436
rect 258350 335424 258356 335436
rect 252244 335396 258356 335424
rect 252244 335384 252250 335396
rect 258350 335384 258356 335396
rect 258408 335384 258414 335436
rect 274818 335384 274824 335436
rect 274876 335424 274882 335436
rect 275002 335424 275008 335436
rect 274876 335396 275008 335424
rect 274876 335384 274882 335396
rect 275002 335384 275008 335396
rect 275060 335384 275066 335436
rect 276106 335384 276112 335436
rect 276164 335424 276170 335436
rect 276658 335424 276664 335436
rect 276164 335396 276664 335424
rect 276164 335384 276170 335396
rect 276658 335384 276664 335396
rect 276716 335384 276722 335436
rect 254486 335316 254492 335368
rect 254544 335356 254550 335368
rect 260834 335356 260840 335368
rect 254544 335328 260840 335356
rect 254544 335316 254550 335328
rect 260834 335316 260840 335328
rect 260892 335316 260898 335368
rect 274726 335316 274732 335368
rect 274784 335356 274790 335368
rect 275370 335356 275376 335368
rect 274784 335328 275376 335356
rect 274784 335316 274790 335328
rect 275370 335316 275376 335328
rect 275428 335316 275434 335368
rect 275830 335316 275836 335368
rect 275888 335356 275894 335368
rect 283742 335356 283748 335368
rect 275888 335328 283748 335356
rect 275888 335316 275894 335328
rect 283742 335316 283748 335328
rect 283800 335316 283806 335368
rect 285674 335316 285680 335368
rect 285732 335356 285738 335368
rect 286410 335356 286416 335368
rect 285732 335328 286416 335356
rect 285732 335316 285738 335328
rect 286410 335316 286416 335328
rect 286468 335316 286474 335368
rect 288342 335316 288348 335368
rect 288400 335356 288406 335368
rect 291838 335356 291844 335368
rect 288400 335328 291844 335356
rect 288400 335316 288406 335328
rect 291838 335316 291844 335328
rect 291896 335316 291902 335368
rect 255682 335248 255688 335300
rect 255740 335288 255746 335300
rect 256326 335288 256332 335300
rect 255740 335260 256332 335288
rect 255740 335248 255746 335260
rect 256326 335248 256332 335260
rect 256384 335248 256390 335300
rect 272334 335248 272340 335300
rect 272392 335288 272398 335300
rect 346854 335288 346860 335300
rect 272392 335260 346860 335288
rect 272392 335248 272398 335260
rect 346854 335248 346860 335260
rect 346912 335248 346918 335300
rect 242894 335180 242900 335232
rect 242952 335220 242958 335232
rect 257890 335220 257896 335232
rect 242952 335192 257896 335220
rect 242952 335180 242958 335192
rect 257890 335180 257896 335192
rect 257948 335180 257954 335232
rect 274266 335180 274272 335232
rect 274324 335220 274330 335232
rect 349154 335220 349160 335232
rect 274324 335192 349160 335220
rect 274324 335180 274330 335192
rect 349154 335180 349160 335192
rect 349212 335180 349218 335232
rect 242250 335112 242256 335164
rect 242308 335152 242314 335164
rect 259914 335152 259920 335164
rect 242308 335124 259920 335152
rect 242308 335112 242314 335124
rect 259914 335112 259920 335124
rect 259972 335112 259978 335164
rect 272702 335112 272708 335164
rect 272760 335152 272766 335164
rect 351914 335152 351920 335164
rect 272760 335124 351920 335152
rect 272760 335112 272766 335124
rect 351914 335112 351920 335124
rect 351972 335112 351978 335164
rect 233234 335044 233240 335096
rect 233292 335084 233298 335096
rect 263410 335084 263416 335096
rect 233292 335056 263416 335084
rect 233292 335044 233298 335056
rect 263410 335044 263416 335056
rect 263468 335044 263474 335096
rect 283466 335044 283472 335096
rect 283524 335084 283530 335096
rect 491294 335084 491300 335096
rect 283524 335056 491300 335084
rect 283524 335044 283530 335056
rect 491294 335044 491300 335056
rect 491352 335044 491358 335096
rect 229094 334976 229100 335028
rect 229152 335016 229158 335028
rect 263042 335016 263048 335028
rect 229152 334988 263048 335016
rect 229152 334976 229158 334988
rect 263042 334976 263048 334988
rect 263100 334976 263106 335028
rect 285582 334976 285588 335028
rect 285640 335016 285646 335028
rect 509234 335016 509240 335028
rect 285640 334988 509240 335016
rect 285640 334976 285646 334988
rect 509234 334976 509240 334988
rect 509292 334976 509298 335028
rect 211154 334908 211160 334960
rect 211212 334948 211218 334960
rect 248966 334948 248972 334960
rect 211212 334920 248972 334948
rect 211212 334908 211218 334920
rect 248966 334908 248972 334920
rect 249024 334908 249030 334960
rect 249242 334908 249248 334960
rect 249300 334948 249306 334960
rect 249426 334948 249432 334960
rect 249300 334920 249432 334948
rect 249300 334908 249306 334920
rect 249426 334908 249432 334920
rect 249484 334908 249490 334960
rect 258810 334948 258816 334960
rect 253906 334920 258816 334948
rect 173894 334840 173900 334892
rect 173952 334880 173958 334892
rect 253906 334880 253934 334920
rect 258810 334908 258816 334920
rect 258868 334908 258874 334960
rect 274542 334908 274548 334960
rect 274600 334948 274606 334960
rect 279878 334948 279884 334960
rect 274600 334920 279884 334948
rect 274600 334908 274606 334920
rect 279878 334908 279884 334920
rect 279936 334908 279942 334960
rect 286226 334908 286232 334960
rect 286284 334948 286290 334960
rect 523034 334948 523040 334960
rect 286284 334920 523040 334948
rect 286284 334908 286290 334920
rect 523034 334908 523040 334920
rect 523092 334908 523098 334960
rect 257154 334880 257160 334892
rect 173952 334852 253934 334880
rect 254642 334852 257160 334880
rect 173952 334840 173958 334852
rect 151814 334772 151820 334824
rect 151872 334812 151878 334824
rect 254642 334812 254670 334852
rect 257154 334840 257160 334852
rect 257212 334840 257218 334892
rect 286686 334840 286692 334892
rect 286744 334880 286750 334892
rect 531314 334880 531320 334892
rect 286744 334852 531320 334880
rect 286744 334840 286750 334852
rect 531314 334840 531320 334852
rect 531372 334840 531378 334892
rect 256050 334812 256056 334824
rect 151872 334784 254670 334812
rect 254734 334784 256056 334812
rect 151872 334772 151878 334784
rect 136634 334704 136640 334756
rect 136692 334744 136698 334756
rect 254734 334744 254762 334784
rect 256050 334772 256056 334784
rect 256108 334772 256114 334824
rect 290918 334772 290924 334824
rect 290976 334812 290982 334824
rect 538214 334812 538220 334824
rect 290976 334784 538220 334812
rect 290976 334772 290982 334784
rect 538214 334772 538220 334784
rect 538272 334772 538278 334824
rect 255958 334744 255964 334756
rect 136692 334716 254762 334744
rect 254826 334716 255964 334744
rect 136692 334704 136698 334716
rect 133874 334636 133880 334688
rect 133932 334676 133938 334688
rect 254826 334676 254854 334716
rect 255958 334704 255964 334716
rect 256016 334704 256022 334756
rect 291010 334704 291016 334756
rect 291068 334744 291074 334756
rect 545114 334744 545120 334756
rect 291068 334716 545120 334744
rect 291068 334704 291074 334716
rect 545114 334704 545120 334716
rect 545172 334704 545178 334756
rect 133932 334648 254854 334676
rect 133932 334636 133938 334648
rect 288618 334636 288624 334688
rect 288676 334676 288682 334688
rect 556154 334676 556160 334688
rect 288676 334648 556160 334676
rect 288676 334636 288682 334648
rect 556154 334636 556160 334648
rect 556212 334636 556218 334688
rect 249242 334568 249248 334620
rect 249300 334608 249306 334620
rect 251358 334608 251364 334620
rect 249300 334580 251364 334608
rect 249300 334568 249306 334580
rect 251358 334568 251364 334580
rect 251416 334568 251422 334620
rect 253198 334568 253204 334620
rect 253256 334608 253262 334620
rect 253474 334608 253480 334620
rect 253256 334580 253480 334608
rect 253256 334568 253262 334580
rect 253474 334568 253480 334580
rect 253532 334568 253538 334620
rect 253934 334568 253940 334620
rect 253992 334608 253998 334620
rect 255130 334608 255136 334620
rect 253992 334580 255136 334608
rect 253992 334568 253998 334580
rect 255130 334568 255136 334580
rect 255188 334568 255194 334620
rect 264238 334568 264244 334620
rect 264296 334608 264302 334620
rect 264606 334608 264612 334620
rect 264296 334580 264612 334608
rect 264296 334568 264302 334580
rect 264606 334568 264612 334580
rect 264664 334568 264670 334620
rect 265434 334568 265440 334620
rect 265492 334608 265498 334620
rect 265802 334608 265808 334620
rect 265492 334580 265808 334608
rect 265492 334568 265498 334580
rect 265802 334568 265808 334580
rect 265860 334568 265866 334620
rect 266722 334568 266728 334620
rect 266780 334608 266786 334620
rect 267182 334608 267188 334620
rect 266780 334580 267188 334608
rect 266780 334568 266786 334580
rect 267182 334568 267188 334580
rect 267240 334568 267246 334620
rect 283190 334568 283196 334620
rect 283248 334608 283254 334620
rect 283374 334608 283380 334620
rect 283248 334580 283380 334608
rect 283248 334568 283254 334580
rect 283374 334568 283380 334580
rect 283432 334568 283438 334620
rect 284386 334568 284392 334620
rect 284444 334608 284450 334620
rect 284846 334608 284852 334620
rect 284444 334580 284852 334608
rect 284444 334568 284450 334580
rect 284846 334568 284852 334580
rect 284904 334568 284910 334620
rect 289630 334568 289636 334620
rect 289688 334608 289694 334620
rect 565814 334608 565820 334620
rect 289688 334580 565820 334608
rect 289688 334568 289694 334580
rect 565814 334568 565820 334580
rect 565872 334568 565878 334620
rect 52454 334500 52460 334552
rect 52512 334540 52518 334552
rect 247034 334540 247040 334552
rect 52512 334512 247040 334540
rect 52512 334500 52518 334512
rect 247034 334500 247040 334512
rect 247092 334500 247098 334552
rect 248874 334500 248880 334552
rect 248932 334540 248938 334552
rect 249150 334540 249156 334552
rect 248932 334512 249156 334540
rect 248932 334500 248938 334512
rect 249150 334500 249156 334512
rect 249208 334500 249214 334552
rect 273806 334432 273812 334484
rect 273864 334472 273870 334484
rect 276750 334472 276756 334484
rect 273864 334444 276756 334472
rect 273864 334432 273870 334444
rect 276750 334432 276756 334444
rect 276808 334432 276814 334484
rect 249150 334364 249156 334416
rect 249208 334404 249214 334416
rect 258994 334404 259000 334416
rect 249208 334376 259000 334404
rect 249208 334364 249214 334376
rect 258994 334364 259000 334376
rect 259052 334364 259058 334416
rect 288526 334364 288532 334416
rect 288584 334404 288590 334416
rect 289354 334404 289360 334416
rect 288584 334376 289360 334404
rect 288584 334364 288590 334376
rect 289354 334364 289360 334376
rect 289412 334364 289418 334416
rect 265710 334228 265716 334280
rect 265768 334268 265774 334280
rect 266262 334268 266268 334280
rect 265768 334240 266268 334268
rect 265768 334228 265774 334240
rect 266262 334228 266268 334240
rect 266320 334228 266326 334280
rect 285766 334024 285772 334076
rect 285824 334064 285830 334076
rect 286594 334064 286600 334076
rect 285824 334036 286600 334064
rect 285824 334024 285830 334036
rect 286594 334024 286600 334036
rect 286652 334024 286658 334076
rect 257264 333900 263594 333928
rect 149054 333820 149060 333872
rect 149112 333860 149118 333872
rect 256694 333860 256700 333872
rect 149112 333832 256700 333860
rect 149112 333820 149118 333832
rect 256694 333820 256700 333832
rect 256752 333820 256758 333872
rect 241514 333752 241520 333804
rect 241572 333792 241578 333804
rect 257264 333792 257292 333900
rect 261202 333792 261208 333804
rect 241572 333764 257292 333792
rect 257356 333764 261208 333792
rect 241572 333752 241578 333764
rect 216674 333684 216680 333736
rect 216732 333724 216738 333736
rect 257356 333724 257384 333764
rect 261202 333752 261208 333764
rect 261260 333752 261266 333804
rect 263566 333792 263594 333900
rect 263962 333792 263968 333804
rect 263566 333764 263968 333792
rect 263962 333752 263968 333764
rect 264020 333752 264026 333804
rect 216732 333696 257384 333724
rect 216732 333684 216738 333696
rect 155954 333616 155960 333668
rect 156012 333656 156018 333668
rect 257522 333656 257528 333668
rect 156012 333628 257528 333656
rect 156012 333616 156018 333628
rect 257522 333616 257528 333628
rect 257580 333616 257586 333668
rect 255314 333548 255320 333600
rect 255372 333588 255378 333600
rect 256418 333588 256424 333600
rect 255372 333560 256424 333588
rect 255372 333548 255378 333560
rect 256418 333548 256424 333560
rect 256476 333548 256482 333600
rect 257430 333548 257436 333600
rect 257488 333588 257494 333600
rect 301130 333588 301136 333600
rect 257488 333560 301136 333588
rect 257488 333548 257494 333560
rect 301130 333548 301136 333560
rect 301188 333548 301194 333600
rect 135254 333480 135260 333532
rect 135312 333520 135318 333532
rect 255590 333520 255596 333532
rect 135312 333492 255596 333520
rect 135312 333480 135318 333492
rect 255590 333480 255596 333492
rect 255648 333480 255654 333532
rect 276474 333480 276480 333532
rect 276532 333520 276538 333532
rect 398834 333520 398840 333532
rect 276532 333492 398840 333520
rect 276532 333480 276538 333492
rect 398834 333480 398840 333492
rect 398892 333480 398898 333532
rect 118694 333412 118700 333464
rect 118752 333452 118758 333464
rect 254578 333452 254584 333464
rect 118752 333424 254584 333452
rect 118752 333412 118758 333424
rect 254578 333412 254584 333424
rect 254636 333412 254642 333464
rect 265618 333452 265624 333464
rect 256252 333424 265624 333452
rect 256252 333396 256280 333424
rect 265618 333412 265624 333424
rect 265676 333412 265682 333464
rect 276934 333412 276940 333464
rect 276992 333452 276998 333464
rect 407114 333452 407120 333464
rect 276992 333424 407120 333452
rect 276992 333412 276998 333424
rect 407114 333412 407120 333424
rect 407172 333412 407178 333464
rect 91094 333344 91100 333396
rect 91152 333384 91158 333396
rect 252278 333384 252284 333396
rect 91152 333356 252284 333384
rect 91152 333344 91158 333356
rect 252278 333344 252284 333356
rect 252336 333344 252342 333396
rect 256234 333344 256240 333396
rect 256292 333344 256298 333396
rect 273806 333344 273812 333396
rect 273864 333384 273870 333396
rect 274174 333384 274180 333396
rect 273864 333356 274180 333384
rect 273864 333344 273870 333356
rect 274174 333344 274180 333356
rect 274232 333344 274238 333396
rect 278958 333344 278964 333396
rect 279016 333384 279022 333396
rect 414014 333384 414020 333396
rect 279016 333356 414020 333384
rect 279016 333344 279022 333356
rect 414014 333344 414020 333356
rect 414072 333344 414078 333396
rect 84194 333276 84200 333328
rect 84252 333316 84258 333328
rect 251542 333316 251548 333328
rect 84252 333288 251548 333316
rect 84252 333276 84258 333288
rect 251542 333276 251548 333288
rect 251600 333276 251606 333328
rect 279142 333276 279148 333328
rect 279200 333316 279206 333328
rect 420914 333316 420920 333328
rect 279200 333288 420920 333316
rect 279200 333276 279206 333288
rect 420914 333276 420920 333288
rect 420972 333276 420978 333328
rect 41414 333208 41420 333260
rect 41472 333248 41478 333260
rect 245378 333248 245384 333260
rect 41472 333220 245384 333248
rect 41472 333208 41478 333220
rect 245378 333208 245384 333220
rect 245436 333208 245442 333260
rect 247126 333208 247132 333260
rect 247184 333248 247190 333260
rect 248046 333248 248052 333260
rect 247184 333220 248052 333248
rect 247184 333208 247190 333220
rect 248046 333208 248052 333220
rect 248104 333208 248110 333260
rect 250070 333208 250076 333260
rect 250128 333248 250134 333260
rect 250254 333248 250260 333260
rect 250128 333220 250260 333248
rect 250128 333208 250134 333220
rect 250254 333208 250260 333220
rect 250312 333208 250318 333260
rect 250346 333208 250352 333260
rect 250404 333248 250410 333260
rect 250714 333248 250720 333260
rect 250404 333220 250720 333248
rect 250404 333208 250410 333220
rect 250714 333208 250720 333220
rect 250772 333208 250778 333260
rect 271966 333208 271972 333260
rect 272024 333248 272030 333260
rect 272242 333248 272248 333260
rect 272024 333220 272248 333248
rect 272024 333208 272030 333220
rect 272242 333208 272248 333220
rect 272300 333208 272306 333260
rect 272518 333208 272524 333260
rect 272576 333248 272582 333260
rect 274174 333248 274180 333260
rect 272576 333220 274180 333248
rect 272576 333208 272582 333220
rect 274174 333208 274180 333220
rect 274232 333208 274238 333260
rect 277578 333208 277584 333260
rect 277636 333248 277642 333260
rect 278314 333248 278320 333260
rect 277636 333220 278320 333248
rect 277636 333208 277642 333220
rect 278314 333208 278320 333220
rect 278372 333208 278378 333260
rect 280062 333208 280068 333260
rect 280120 333248 280126 333260
rect 438854 333248 438860 333260
rect 280120 333220 438860 333248
rect 280120 333208 280126 333220
rect 438854 333208 438860 333220
rect 438912 333208 438918 333260
rect 247770 333140 247776 333192
rect 247828 333180 247834 333192
rect 248782 333180 248788 333192
rect 247828 333152 248788 333180
rect 247828 333140 247834 333152
rect 248782 333140 248788 333152
rect 248840 333140 248846 333192
rect 249978 333140 249984 333192
rect 250036 333180 250042 333192
rect 250806 333180 250812 333192
rect 250036 333152 250812 333180
rect 250036 333140 250042 333152
rect 250806 333140 250812 333152
rect 250864 333140 250870 333192
rect 274358 333140 274364 333192
rect 274416 333180 274422 333192
rect 276566 333180 276572 333192
rect 274416 333152 276572 333180
rect 274416 333140 274422 333152
rect 276566 333140 276572 333152
rect 276624 333140 276630 333192
rect 248690 333072 248696 333124
rect 248748 333112 248754 333124
rect 249426 333112 249432 333124
rect 248748 333084 249432 333112
rect 248748 333072 248754 333084
rect 249426 333072 249432 333084
rect 249484 333072 249490 333124
rect 250254 333072 250260 333124
rect 250312 333112 250318 333124
rect 250990 333112 250996 333124
rect 250312 333084 250996 333112
rect 250312 333072 250318 333084
rect 250990 333072 250996 333084
rect 251048 333072 251054 333124
rect 247402 333004 247408 333056
rect 247460 333044 247466 333056
rect 247954 333044 247960 333056
rect 247460 333016 247960 333044
rect 247460 333004 247466 333016
rect 247954 333004 247960 333016
rect 248012 333004 248018 333056
rect 248782 333004 248788 333056
rect 248840 333044 248846 333056
rect 249610 333044 249616 333056
rect 248840 333016 249616 333044
rect 248840 333004 248846 333016
rect 249610 333004 249616 333016
rect 249668 333004 249674 333056
rect 272426 333004 272432 333056
rect 272484 333044 272490 333056
rect 272610 333044 272616 333056
rect 272484 333016 272616 333044
rect 272484 333004 272490 333016
rect 272610 333004 272616 333016
rect 272668 333004 272674 333056
rect 246758 332936 246764 332988
rect 246816 332976 246822 332988
rect 265802 332976 265808 332988
rect 246816 332948 265808 332976
rect 246816 332936 246822 332948
rect 265802 332936 265808 332948
rect 265860 332936 265866 332988
rect 273530 332868 273536 332920
rect 273588 332908 273594 332920
rect 274082 332908 274088 332920
rect 273588 332880 274088 332908
rect 273588 332868 273594 332880
rect 274082 332868 274088 332880
rect 274140 332868 274146 332920
rect 243630 332324 243636 332376
rect 243688 332364 243694 332376
rect 260742 332364 260748 332376
rect 243688 332336 260748 332364
rect 243688 332324 243694 332336
rect 260742 332324 260748 332336
rect 260800 332324 260806 332376
rect 226334 332256 226340 332308
rect 226392 332296 226398 332308
rect 262674 332296 262680 332308
rect 226392 332268 262680 332296
rect 226392 332256 226398 332268
rect 262674 332256 262680 332268
rect 262732 332256 262738 332308
rect 233878 332188 233884 332240
rect 233936 332228 233942 332240
rect 258534 332228 258540 332240
rect 233936 332200 258540 332228
rect 233936 332188 233942 332200
rect 258534 332188 258540 332200
rect 258592 332188 258598 332240
rect 259914 332188 259920 332240
rect 259972 332228 259978 332240
rect 300946 332228 300952 332240
rect 259972 332200 300952 332228
rect 259972 332188 259978 332200
rect 300946 332188 300952 332200
rect 301004 332188 301010 332240
rect 257798 332120 257804 332172
rect 257856 332160 257862 332172
rect 301038 332160 301044 332172
rect 257856 332132 301044 332160
rect 257856 332120 257862 332132
rect 301038 332120 301044 332132
rect 301096 332120 301102 332172
rect 168374 332052 168380 332104
rect 168432 332092 168438 332104
rect 246850 332092 246856 332104
rect 168432 332064 246856 332092
rect 168432 332052 168438 332064
rect 246850 332052 246856 332064
rect 246908 332052 246914 332104
rect 272978 332052 272984 332104
rect 273036 332092 273042 332104
rect 354674 332092 354680 332104
rect 273036 332064 354680 332092
rect 273036 332052 273042 332064
rect 354674 332052 354680 332064
rect 354732 332052 354738 332104
rect 122834 331984 122840 332036
rect 122892 332024 122898 332036
rect 255406 332024 255412 332036
rect 122892 331996 255412 332024
rect 122892 331984 122898 331996
rect 255406 331984 255412 331996
rect 255464 331984 255470 332036
rect 281810 331984 281816 332036
rect 281868 332024 281874 332036
rect 379514 332024 379520 332036
rect 281868 331996 379520 332024
rect 281868 331984 281874 331996
rect 379514 331984 379520 331996
rect 379572 331984 379578 332036
rect 74534 331916 74540 331968
rect 74592 331956 74598 331968
rect 251174 331956 251180 331968
rect 74592 331928 251180 331956
rect 74592 331916 74598 331928
rect 251174 331916 251180 331928
rect 251232 331916 251238 331968
rect 289078 331916 289084 331968
rect 289136 331956 289142 331968
rect 556246 331956 556252 331968
rect 289136 331928 556252 331956
rect 289136 331916 289142 331928
rect 556246 331916 556252 331928
rect 556304 331916 556310 331968
rect 34514 331848 34520 331900
rect 34572 331888 34578 331900
rect 247586 331888 247592 331900
rect 34572 331860 247592 331888
rect 34572 331848 34578 331860
rect 247586 331848 247592 331860
rect 247644 331848 247650 331900
rect 289170 331848 289176 331900
rect 289228 331888 289234 331900
rect 564434 331888 564440 331900
rect 289228 331860 564440 331888
rect 289228 331848 289234 331860
rect 564434 331848 564440 331860
rect 564492 331848 564498 331900
rect 248966 331644 248972 331696
rect 249024 331684 249030 331696
rect 249702 331684 249708 331696
rect 249024 331656 249708 331684
rect 249024 331644 249030 331656
rect 249702 331644 249708 331656
rect 249760 331644 249766 331696
rect 260742 331236 260748 331288
rect 260800 331276 260806 331288
rect 265986 331276 265992 331288
rect 260800 331248 265992 331276
rect 260800 331236 260806 331248
rect 265986 331236 265992 331248
rect 266044 331236 266050 331288
rect 257246 331168 257252 331220
rect 257304 331208 257310 331220
rect 257522 331208 257528 331220
rect 257304 331180 257528 331208
rect 257304 331168 257310 331180
rect 257522 331168 257528 331180
rect 257580 331168 257586 331220
rect 251634 330964 251640 331016
rect 251692 331004 251698 331016
rect 251910 331004 251916 331016
rect 251692 330976 251916 331004
rect 251692 330964 251698 330976
rect 251910 330964 251916 330976
rect 251968 330964 251974 331016
rect 272150 330964 272156 331016
rect 272208 331004 272214 331016
rect 272794 331004 272800 331016
rect 272208 330976 272800 331004
rect 272208 330964 272214 330976
rect 272794 330964 272800 330976
rect 272852 330964 272858 331016
rect 251174 330896 251180 330948
rect 251232 330936 251238 330948
rect 252462 330936 252468 330948
rect 251232 330908 252468 330936
rect 251232 330896 251238 330908
rect 252462 330896 252468 330908
rect 252520 330896 252526 330948
rect 234706 330828 234712 330880
rect 234764 330868 234770 330880
rect 263410 330868 263416 330880
rect 234764 330840 263416 330868
rect 234764 330828 234770 330840
rect 263410 330828 263416 330840
rect 263468 330828 263474 330880
rect 207014 330760 207020 330812
rect 207072 330800 207078 330812
rect 261294 330800 261300 330812
rect 207072 330772 261300 330800
rect 207072 330760 207078 330772
rect 261294 330760 261300 330772
rect 261352 330760 261358 330812
rect 266446 330760 266452 330812
rect 266504 330760 266510 330812
rect 269114 330760 269120 330812
rect 269172 330800 269178 330812
rect 270218 330800 270224 330812
rect 269172 330772 270224 330800
rect 269172 330760 269178 330772
rect 270218 330760 270224 330772
rect 270276 330760 270282 330812
rect 193214 330692 193220 330744
rect 193272 330732 193278 330744
rect 259546 330732 259552 330744
rect 193272 330704 259552 330732
rect 193272 330692 193278 330704
rect 259546 330692 259552 330704
rect 259604 330692 259610 330744
rect 264882 330732 264888 330744
rect 263566 330704 264888 330732
rect 184934 330624 184940 330676
rect 184992 330664 184998 330676
rect 251174 330664 251180 330676
rect 184992 330636 251180 330664
rect 184992 330624 184998 330636
rect 251174 330624 251180 330636
rect 251232 330624 251238 330676
rect 251358 330624 251364 330676
rect 251416 330664 251422 330676
rect 252002 330664 252008 330676
rect 251416 330636 252008 330664
rect 251416 330624 251422 330636
rect 252002 330624 252008 330636
rect 252060 330624 252066 330676
rect 252830 330624 252836 330676
rect 252888 330664 252894 330676
rect 253106 330664 253112 330676
rect 252888 330636 253112 330664
rect 252888 330624 252894 330636
rect 253106 330624 253112 330636
rect 253164 330624 253170 330676
rect 255958 330624 255964 330676
rect 256016 330664 256022 330676
rect 263566 330664 263594 330704
rect 264882 330692 264888 330704
rect 264940 330692 264946 330744
rect 256016 330636 263594 330664
rect 256016 330624 256022 330636
rect 263778 330624 263784 330676
rect 263836 330664 263842 330676
rect 264330 330664 264336 330676
rect 263836 330636 264336 330664
rect 263836 330624 263842 330636
rect 264330 330624 264336 330636
rect 264388 330624 264394 330676
rect 189074 330556 189080 330608
rect 189132 330596 189138 330608
rect 260282 330596 260288 330608
rect 189132 330568 260288 330596
rect 189132 330556 189138 330568
rect 260282 330556 260288 330568
rect 260340 330556 260346 330608
rect 263962 330556 263968 330608
rect 264020 330596 264026 330608
rect 264790 330596 264796 330608
rect 264020 330568 264796 330596
rect 264020 330556 264026 330568
rect 264790 330556 264796 330568
rect 264848 330556 264854 330608
rect 266464 330596 266492 330760
rect 269298 330692 269304 330744
rect 269356 330732 269362 330744
rect 270034 330732 270040 330744
rect 269356 330704 270040 330732
rect 269356 330692 269362 330704
rect 270034 330692 270040 330704
rect 270092 330692 270098 330744
rect 266906 330624 266912 330676
rect 266964 330664 266970 330676
rect 266964 330636 267044 330664
rect 266964 330624 266970 330636
rect 266538 330596 266544 330608
rect 266464 330568 266544 330596
rect 266538 330556 266544 330568
rect 266596 330556 266602 330608
rect 60734 330488 60740 330540
rect 60792 330528 60798 330540
rect 245746 330528 245752 330540
rect 60792 330500 245752 330528
rect 60792 330488 60798 330500
rect 245746 330488 245752 330500
rect 245804 330488 245810 330540
rect 245838 330488 245844 330540
rect 245896 330528 245902 330540
rect 246574 330528 246580 330540
rect 245896 330500 246580 330528
rect 245896 330488 245902 330500
rect 246574 330488 246580 330500
rect 246632 330488 246638 330540
rect 247862 330488 247868 330540
rect 247920 330528 247926 330540
rect 248322 330528 248328 330540
rect 247920 330500 248328 330528
rect 247920 330488 247926 330500
rect 248322 330488 248328 330500
rect 248380 330488 248386 330540
rect 251542 330488 251548 330540
rect 251600 330528 251606 330540
rect 252094 330528 252100 330540
rect 251600 330500 252100 330528
rect 251600 330488 251606 330500
rect 252094 330488 252100 330500
rect 252152 330488 252158 330540
rect 252554 330488 252560 330540
rect 252612 330528 252618 330540
rect 252830 330528 252836 330540
rect 252612 330500 252836 330528
rect 252612 330488 252618 330500
rect 252830 330488 252836 330500
rect 252888 330488 252894 330540
rect 253290 330488 253296 330540
rect 253348 330528 253354 330540
rect 253750 330528 253756 330540
rect 253348 330500 253756 330528
rect 253348 330488 253354 330500
rect 253750 330488 253756 330500
rect 253808 330488 253814 330540
rect 264054 330488 264060 330540
rect 264112 330528 264118 330540
rect 264330 330528 264336 330540
rect 264112 330500 264336 330528
rect 264112 330488 264118 330500
rect 264330 330488 264336 330500
rect 264388 330488 264394 330540
rect 265250 330488 265256 330540
rect 265308 330528 265314 330540
rect 265526 330528 265532 330540
rect 265308 330500 265532 330528
rect 265308 330488 265314 330500
rect 265526 330488 265532 330500
rect 265584 330488 265590 330540
rect 267016 330472 267044 330636
rect 269114 330624 269120 330676
rect 269172 330664 269178 330676
rect 269574 330664 269580 330676
rect 269172 330636 269580 330664
rect 269172 330624 269178 330636
rect 269574 330624 269580 330636
rect 269632 330624 269638 330676
rect 271138 330664 271144 330676
rect 271064 330636 271144 330664
rect 268286 330488 268292 330540
rect 268344 330528 268350 330540
rect 268470 330528 268476 330540
rect 268344 330500 268476 330528
rect 268344 330488 268350 330500
rect 268470 330488 268476 330500
rect 268528 330488 268534 330540
rect 269574 330488 269580 330540
rect 269632 330528 269638 330540
rect 269850 330528 269856 330540
rect 269632 330500 269856 330528
rect 269632 330488 269638 330500
rect 269850 330488 269856 330500
rect 269908 330488 269914 330540
rect 271064 330472 271092 330636
rect 271138 330624 271144 330636
rect 271196 330624 271202 330676
rect 281350 330624 281356 330676
rect 281408 330664 281414 330676
rect 361574 330664 361580 330676
rect 281408 330636 361580 330664
rect 281408 330624 281414 330636
rect 361574 330624 361580 330636
rect 361632 330624 361638 330676
rect 275646 330556 275652 330608
rect 275704 330596 275710 330608
rect 358814 330596 358820 330608
rect 275704 330568 358820 330596
rect 275704 330556 275710 330568
rect 358814 330556 358820 330568
rect 358872 330556 358878 330608
rect 290826 330488 290832 330540
rect 290884 330528 290890 330540
rect 572714 330528 572720 330540
rect 290884 330500 572720 330528
rect 290884 330488 290890 330500
rect 572714 330488 572720 330500
rect 572772 330488 572778 330540
rect 246114 330420 246120 330472
rect 246172 330460 246178 330472
rect 246666 330460 246672 330472
rect 246172 330432 246672 330460
rect 246172 330420 246178 330432
rect 246666 330420 246672 330432
rect 246724 330420 246730 330472
rect 251450 330420 251456 330472
rect 251508 330460 251514 330472
rect 252370 330460 252376 330472
rect 251508 330432 252376 330460
rect 251508 330420 251514 330432
rect 252370 330420 252376 330432
rect 252428 330420 252434 330472
rect 253014 330420 253020 330472
rect 253072 330460 253078 330472
rect 253842 330460 253848 330472
rect 253072 330432 253848 330460
rect 253072 330420 253078 330432
rect 253842 330420 253848 330432
rect 253900 330420 253906 330472
rect 263870 330420 263876 330472
rect 263928 330460 263934 330472
rect 264422 330460 264428 330472
rect 263928 330432 264428 330460
rect 263928 330420 263934 330432
rect 264422 330420 264428 330432
rect 264480 330420 264486 330472
rect 266998 330420 267004 330472
rect 267056 330420 267062 330472
rect 268010 330420 268016 330472
rect 268068 330460 268074 330472
rect 268194 330460 268200 330472
rect 268068 330432 268200 330460
rect 268068 330420 268074 330432
rect 268194 330420 268200 330432
rect 268252 330420 268258 330472
rect 269206 330420 269212 330472
rect 269264 330460 269270 330472
rect 269390 330460 269396 330472
rect 269264 330432 269396 330460
rect 269264 330420 269270 330432
rect 269390 330420 269396 330432
rect 269448 330420 269454 330472
rect 269482 330420 269488 330472
rect 269540 330460 269546 330472
rect 269942 330460 269948 330472
rect 269540 330432 269948 330460
rect 269540 330420 269546 330432
rect 269942 330420 269948 330432
rect 270000 330420 270006 330472
rect 271046 330420 271052 330472
rect 271104 330420 271110 330472
rect 245746 330352 245752 330404
rect 245804 330392 245810 330404
rect 246942 330392 246948 330404
rect 245804 330364 246948 330392
rect 245804 330352 245810 330364
rect 246942 330352 246948 330364
rect 247000 330352 247006 330404
rect 252646 330352 252652 330404
rect 252704 330392 252710 330404
rect 253658 330392 253664 330404
rect 252704 330364 253664 330392
rect 252704 330352 252710 330364
rect 253658 330352 253664 330364
rect 253716 330352 253722 330404
rect 264054 330352 264060 330404
rect 264112 330392 264118 330404
rect 264514 330392 264520 330404
rect 264112 330364 264520 330392
rect 264112 330352 264118 330364
rect 264514 330352 264520 330364
rect 264572 330352 264578 330404
rect 265526 330352 265532 330404
rect 265584 330392 265590 330404
rect 266078 330392 266084 330404
rect 265584 330364 266084 330392
rect 265584 330352 265590 330364
rect 266078 330352 266084 330364
rect 266136 330352 266142 330404
rect 266722 330352 266728 330404
rect 266780 330392 266786 330404
rect 267366 330392 267372 330404
rect 266780 330364 267372 330392
rect 266780 330352 266786 330364
rect 267366 330352 267372 330364
rect 267424 330352 267430 330404
rect 268286 330352 268292 330404
rect 268344 330392 268350 330404
rect 268562 330392 268568 330404
rect 268344 330364 268568 330392
rect 268344 330352 268350 330364
rect 268562 330352 268568 330364
rect 268620 330352 268626 330404
rect 270862 330352 270868 330404
rect 270920 330392 270926 330404
rect 271322 330392 271328 330404
rect 270920 330364 271328 330392
rect 270920 330352 270926 330364
rect 271322 330352 271328 330364
rect 271380 330352 271386 330404
rect 251634 330284 251640 330336
rect 251692 330324 251698 330336
rect 251818 330324 251824 330336
rect 251692 330296 251824 330324
rect 251692 330284 251698 330296
rect 251818 330284 251824 330296
rect 251876 330284 251882 330336
rect 254946 330284 254952 330336
rect 255004 330324 255010 330336
rect 264606 330324 264612 330336
rect 255004 330296 264612 330324
rect 255004 330284 255010 330296
rect 264606 330284 264612 330296
rect 264664 330284 264670 330336
rect 268194 330284 268200 330336
rect 268252 330324 268258 330336
rect 268746 330324 268752 330336
rect 268252 330296 268752 330324
rect 268252 330284 268258 330296
rect 268746 330284 268752 330296
rect 268804 330284 268810 330336
rect 269390 330284 269396 330336
rect 269448 330324 269454 330336
rect 270126 330324 270132 330336
rect 269448 330296 270132 330324
rect 269448 330284 269454 330296
rect 270126 330284 270132 330296
rect 270184 330284 270190 330336
rect 270678 330284 270684 330336
rect 270736 330324 270742 330336
rect 271598 330324 271604 330336
rect 270736 330296 271604 330324
rect 270736 330284 270742 330296
rect 271598 330284 271604 330296
rect 271656 330284 271662 330336
rect 267734 330216 267740 330268
rect 267792 330256 267798 330268
rect 268562 330256 268568 330268
rect 267792 330228 268568 330256
rect 267792 330216 267798 330228
rect 268562 330216 268568 330228
rect 268620 330216 268626 330268
rect 265342 329672 265348 329724
rect 265400 329712 265406 329724
rect 266170 329712 266176 329724
rect 265400 329684 266176 329712
rect 265400 329672 265406 329684
rect 266170 329672 266176 329684
rect 266228 329672 266234 329724
rect 220814 329332 220820 329384
rect 220872 329372 220878 329384
rect 253474 329372 253480 329384
rect 220872 329344 253480 329372
rect 220872 329332 220878 329344
rect 253474 329332 253480 329344
rect 253532 329332 253538 329384
rect 153194 329264 153200 329316
rect 153252 329304 153258 329316
rect 256970 329304 256976 329316
rect 153252 329276 256976 329304
rect 153252 329264 153258 329276
rect 256970 329264 256976 329276
rect 257028 329264 257034 329316
rect 126974 329196 126980 329248
rect 127032 329236 127038 329248
rect 253934 329236 253940 329248
rect 127032 329208 253940 329236
rect 127032 329196 127038 329208
rect 253934 329196 253940 329208
rect 253992 329196 253998 329248
rect 52546 329128 52552 329180
rect 52604 329168 52610 329180
rect 248138 329168 248144 329180
rect 52604 329140 248144 329168
rect 52604 329128 52610 329140
rect 248138 329128 248144 329140
rect 248196 329128 248202 329180
rect 283650 329128 283656 329180
rect 283708 329168 283714 329180
rect 489914 329168 489920 329180
rect 283708 329140 489920 329168
rect 283708 329128 283714 329140
rect 489914 329128 489920 329140
rect 489972 329128 489978 329180
rect 37274 329060 37280 329112
rect 37332 329100 37338 329112
rect 248230 329100 248236 329112
rect 37332 329072 248236 329100
rect 37332 329060 37338 329072
rect 248230 329060 248236 329072
rect 248288 329060 248294 329112
rect 287606 329060 287612 329112
rect 287664 329100 287670 329112
rect 539594 329100 539600 329112
rect 287664 329072 539600 329100
rect 287664 329060 287670 329072
rect 539594 329060 539600 329072
rect 539652 329060 539658 329112
rect 283006 328380 283012 328432
rect 283064 328420 283070 328432
rect 283466 328420 283472 328432
rect 283064 328392 283472 328420
rect 283064 328380 283070 328392
rect 283466 328380 283472 328392
rect 283524 328380 283530 328432
rect 274634 328108 274640 328160
rect 274692 328148 274698 328160
rect 275646 328148 275652 328160
rect 274692 328120 275652 328148
rect 274692 328108 274698 328120
rect 275646 328108 275652 328120
rect 275704 328108 275710 328160
rect 180794 327836 180800 327888
rect 180852 327876 180858 327888
rect 259362 327876 259368 327888
rect 180852 327848 259368 327876
rect 180852 327836 180858 327848
rect 259362 327836 259368 327848
rect 259420 327836 259426 327888
rect 276934 327836 276940 327888
rect 276992 327876 276998 327888
rect 398926 327876 398932 327888
rect 276992 327848 398932 327876
rect 276992 327836 276998 327848
rect 398926 327836 398932 327848
rect 398984 327836 398990 327888
rect 171134 327768 171140 327820
rect 171192 327808 171198 327820
rect 252186 327808 252192 327820
rect 171192 327780 252192 327808
rect 171192 327768 171198 327780
rect 252186 327768 252192 327780
rect 252244 327768 252250 327820
rect 278222 327768 278228 327820
rect 278280 327808 278286 327820
rect 423674 327808 423680 327820
rect 278280 327780 423680 327808
rect 278280 327768 278286 327780
rect 423674 327768 423680 327780
rect 423732 327768 423738 327820
rect 46934 327700 46940 327752
rect 46992 327740 46998 327752
rect 249058 327740 249064 327752
rect 46992 327712 249064 327740
rect 46992 327700 46998 327712
rect 249058 327700 249064 327712
rect 249116 327700 249122 327752
rect 290182 327700 290188 327752
rect 290240 327740 290246 327752
rect 575474 327740 575480 327752
rect 290240 327712 575480 327740
rect 290240 327700 290246 327712
rect 575474 327700 575480 327712
rect 575532 327700 575538 327752
rect 276290 327360 276296 327412
rect 276348 327400 276354 327412
rect 276934 327400 276940 327412
rect 276348 327372 276940 327400
rect 276348 327360 276354 327372
rect 276934 327360 276940 327372
rect 276992 327360 276998 327412
rect 285122 326748 285128 326800
rect 285180 326788 285186 326800
rect 294506 326788 294512 326800
rect 285180 326760 294512 326788
rect 285180 326748 285186 326760
rect 294506 326748 294512 326760
rect 294564 326748 294570 326800
rect 257154 326680 257160 326732
rect 257212 326720 257218 326732
rect 257982 326720 257988 326732
rect 257212 326692 257988 326720
rect 257212 326680 257218 326692
rect 257982 326680 257988 326692
rect 258040 326680 258046 326732
rect 274726 326680 274732 326732
rect 274784 326680 274790 326732
rect 284294 326680 284300 326732
rect 284352 326720 284358 326732
rect 285306 326720 285312 326732
rect 284352 326692 285312 326720
rect 284352 326680 284358 326692
rect 285306 326680 285312 326692
rect 285364 326680 285370 326732
rect 287716 326692 289814 326720
rect 257614 326544 257620 326596
rect 257672 326584 257678 326596
rect 257982 326584 257988 326596
rect 257672 326556 257988 326584
rect 257672 326544 257678 326556
rect 257982 326544 257988 326556
rect 258040 326544 258046 326596
rect 261386 326544 261392 326596
rect 261444 326584 261450 326596
rect 261754 326584 261760 326596
rect 261444 326556 261760 326584
rect 261444 326544 261450 326556
rect 261754 326544 261760 326556
rect 261812 326544 261818 326596
rect 261938 326516 261944 326528
rect 253906 326488 261944 326516
rect 209774 326340 209780 326392
rect 209832 326380 209838 326392
rect 253906 326380 253934 326488
rect 261938 326476 261944 326488
rect 261996 326476 262002 326528
rect 274744 326460 274772 326680
rect 279878 326612 279884 326664
rect 279936 326652 279942 326664
rect 287716 326652 287744 326692
rect 279936 326624 287744 326652
rect 279936 326612 279942 326624
rect 288618 326612 288624 326664
rect 288676 326652 288682 326664
rect 288802 326652 288808 326664
rect 288676 326624 288808 326652
rect 288676 326612 288682 326624
rect 288802 326612 288808 326624
rect 288860 326612 288866 326664
rect 289786 326652 289814 326692
rect 365714 326652 365720 326664
rect 289786 326624 365720 326652
rect 365714 326612 365720 326624
rect 365772 326612 365778 326664
rect 275278 326544 275284 326596
rect 275336 326544 275342 326596
rect 286042 326544 286048 326596
rect 286100 326584 286106 326596
rect 286100 326556 290136 326584
rect 286100 326544 286106 326556
rect 254302 326408 254308 326460
rect 254360 326448 254366 326460
rect 254762 326448 254768 326460
rect 254360 326420 254768 326448
rect 254360 326408 254366 326420
rect 254762 326408 254768 326420
rect 254820 326408 254826 326460
rect 256142 326408 256148 326460
rect 256200 326448 256206 326460
rect 256510 326448 256516 326460
rect 256200 326420 256516 326448
rect 256200 326408 256206 326420
rect 256510 326408 256516 326420
rect 256568 326408 256574 326460
rect 262490 326408 262496 326460
rect 262548 326448 262554 326460
rect 263226 326448 263232 326460
rect 262548 326420 263232 326448
rect 262548 326408 262554 326420
rect 263226 326408 263232 326420
rect 263284 326408 263290 326460
rect 274726 326408 274732 326460
rect 274784 326408 274790 326460
rect 209832 326352 253934 326380
rect 209832 326340 209838 326352
rect 254486 326340 254492 326392
rect 254544 326380 254550 326392
rect 255222 326380 255228 326392
rect 254544 326352 255228 326380
rect 254544 326340 254550 326352
rect 255222 326340 255228 326352
rect 255280 326340 255286 326392
rect 256970 326340 256976 326392
rect 257028 326380 257034 326392
rect 257706 326380 257712 326392
rect 257028 326352 257712 326380
rect 257028 326340 257034 326352
rect 257706 326340 257712 326352
rect 257764 326340 257770 326392
rect 258258 326340 258264 326392
rect 258316 326380 258322 326392
rect 259270 326380 259276 326392
rect 258316 326352 259276 326380
rect 258316 326340 258322 326352
rect 259270 326340 259276 326352
rect 259328 326340 259334 326392
rect 260006 326340 260012 326392
rect 260064 326380 260070 326392
rect 260650 326380 260656 326392
rect 260064 326352 260656 326380
rect 260064 326340 260070 326352
rect 260650 326340 260656 326352
rect 260708 326340 260714 326392
rect 261294 326340 261300 326392
rect 261352 326380 261358 326392
rect 261846 326380 261852 326392
rect 261352 326352 261852 326380
rect 261352 326340 261358 326352
rect 261846 326340 261852 326352
rect 261904 326340 261910 326392
rect 262674 326340 262680 326392
rect 262732 326380 262738 326392
rect 263318 326380 263324 326392
rect 262732 326352 263324 326380
rect 262732 326340 262738 326352
rect 263318 326340 263324 326352
rect 263376 326340 263382 326392
rect 275186 326340 275192 326392
rect 275244 326380 275250 326392
rect 275296 326380 275324 326544
rect 286410 326476 286416 326528
rect 286468 326516 286474 326528
rect 290108 326516 290136 326556
rect 294506 326544 294512 326596
rect 294564 326584 294570 326596
rect 511994 326584 512000 326596
rect 294564 326556 512000 326584
rect 294564 326544 294570 326556
rect 511994 326544 512000 326556
rect 512052 326544 512058 326596
rect 523126 326516 523132 326528
rect 286468 326488 290044 326516
rect 290108 326488 523132 326516
rect 286468 326476 286474 326488
rect 277578 326408 277584 326460
rect 277636 326408 277642 326460
rect 277670 326408 277676 326460
rect 277728 326448 277734 326460
rect 277854 326448 277860 326460
rect 277728 326420 277860 326448
rect 277728 326408 277734 326420
rect 277854 326408 277860 326420
rect 277912 326408 277918 326460
rect 281994 326408 282000 326460
rect 282052 326448 282058 326460
rect 282270 326448 282276 326460
rect 282052 326420 282276 326448
rect 282052 326408 282058 326420
rect 282270 326408 282276 326420
rect 282328 326408 282334 326460
rect 284478 326408 284484 326460
rect 284536 326448 284542 326460
rect 284846 326448 284852 326460
rect 284536 326420 284852 326448
rect 284536 326408 284542 326420
rect 284846 326408 284852 326420
rect 284904 326408 284910 326460
rect 289906 326408 289912 326460
rect 289964 326408 289970 326460
rect 290016 326448 290044 326488
rect 523126 326476 523132 326488
rect 523184 326476 523190 326528
rect 528554 326448 528560 326460
rect 290016 326420 528560 326448
rect 528554 326408 528560 326420
rect 528612 326408 528618 326460
rect 275244 326352 275324 326380
rect 275244 326340 275250 326352
rect 276014 326340 276020 326392
rect 276072 326380 276078 326392
rect 276842 326380 276848 326392
rect 276072 326352 276848 326380
rect 276072 326340 276078 326352
rect 276842 326340 276848 326352
rect 276900 326340 276906 326392
rect 277596 326380 277624 326408
rect 277596 326352 277808 326380
rect 254210 326272 254216 326324
rect 254268 326312 254274 326324
rect 254854 326312 254860 326324
rect 254268 326284 254860 326312
rect 254268 326272 254274 326284
rect 254854 326272 254860 326284
rect 254912 326272 254918 326324
rect 261386 326272 261392 326324
rect 261444 326312 261450 326324
rect 262030 326312 262036 326324
rect 261444 326284 262036 326312
rect 261444 326272 261450 326284
rect 262030 326272 262036 326284
rect 262088 326272 262094 326324
rect 277780 326256 277808 326352
rect 278958 326340 278964 326392
rect 279016 326380 279022 326392
rect 279602 326380 279608 326392
rect 279016 326352 279608 326380
rect 279016 326340 279022 326352
rect 279602 326340 279608 326352
rect 279660 326340 279666 326392
rect 280522 326340 280528 326392
rect 280580 326380 280586 326392
rect 281258 326380 281264 326392
rect 280580 326352 281264 326380
rect 280580 326340 280586 326352
rect 281258 326340 281264 326352
rect 281316 326340 281322 326392
rect 287238 326340 287244 326392
rect 287296 326380 287302 326392
rect 287422 326380 287428 326392
rect 287296 326352 287428 326380
rect 287296 326340 287302 326352
rect 287422 326340 287428 326352
rect 287480 326340 287486 326392
rect 288802 326340 288808 326392
rect 288860 326380 288866 326392
rect 289446 326380 289452 326392
rect 288860 326352 289452 326380
rect 288860 326340 288866 326352
rect 289446 326340 289452 326352
rect 289504 326340 289510 326392
rect 289924 326380 289952 326408
rect 572806 326380 572812 326392
rect 289924 326352 572812 326380
rect 572806 326340 572812 326352
rect 572864 326340 572870 326392
rect 280614 326272 280620 326324
rect 280672 326312 280678 326324
rect 280798 326312 280804 326324
rect 280672 326284 280804 326312
rect 280672 326272 280678 326284
rect 280798 326272 280804 326284
rect 280856 326272 280862 326324
rect 256326 326204 256332 326256
rect 256384 326204 256390 326256
rect 260190 326204 260196 326256
rect 260248 326244 260254 326256
rect 260374 326244 260380 326256
rect 260248 326216 260380 326244
rect 260248 326204 260254 326216
rect 260374 326204 260380 326216
rect 260432 326204 260438 326256
rect 275278 326204 275284 326256
rect 275336 326244 275342 326256
rect 275554 326244 275560 326256
rect 275336 326216 275560 326244
rect 275336 326204 275342 326216
rect 275554 326204 275560 326216
rect 275612 326204 275618 326256
rect 276290 326204 276296 326256
rect 276348 326244 276354 326256
rect 276658 326244 276664 326256
rect 276348 326216 276664 326244
rect 276348 326204 276354 326216
rect 276658 326204 276664 326216
rect 276716 326204 276722 326256
rect 277762 326204 277768 326256
rect 277820 326204 277826 326256
rect 284570 326204 284576 326256
rect 284628 326244 284634 326256
rect 284754 326244 284760 326256
rect 284628 326216 284760 326244
rect 284628 326204 284634 326216
rect 284754 326204 284760 326216
rect 284812 326204 284818 326256
rect 285950 326204 285956 326256
rect 286008 326244 286014 326256
rect 286134 326244 286140 326256
rect 286008 326216 286140 326244
rect 286008 326204 286014 326216
rect 286134 326204 286140 326216
rect 286192 326204 286198 326256
rect 287422 326204 287428 326256
rect 287480 326244 287486 326256
rect 287790 326244 287796 326256
rect 287480 326216 287796 326244
rect 287480 326204 287486 326216
rect 287790 326204 287796 326216
rect 287848 326204 287854 326256
rect 289814 326204 289820 326256
rect 289872 326244 289878 326256
rect 290734 326244 290740 326256
rect 289872 326216 290740 326244
rect 289872 326204 289878 326216
rect 290734 326204 290740 326216
rect 290792 326204 290798 326256
rect 254670 325932 254676 325984
rect 254728 325972 254734 325984
rect 254946 325972 254952 325984
rect 254728 325944 254952 325972
rect 254728 325932 254734 325944
rect 254946 325932 254952 325944
rect 255004 325932 255010 325984
rect 256344 325972 256372 326204
rect 258442 326136 258448 326188
rect 258500 326176 258506 326188
rect 258994 326176 259000 326188
rect 258500 326148 259000 326176
rect 258500 326136 258506 326148
rect 258994 326136 259000 326148
rect 259052 326136 259058 326188
rect 274910 326136 274916 326188
rect 274968 326176 274974 326188
rect 275462 326176 275468 326188
rect 274968 326148 275468 326176
rect 274968 326136 274974 326148
rect 275462 326136 275468 326148
rect 275520 326136 275526 326188
rect 277486 326136 277492 326188
rect 277544 326176 277550 326188
rect 278130 326176 278136 326188
rect 277544 326148 278136 326176
rect 277544 326136 277550 326148
rect 278130 326136 278136 326148
rect 278188 326136 278194 326188
rect 275002 326068 275008 326120
rect 275060 326108 275066 326120
rect 275830 326108 275836 326120
rect 275060 326080 275836 326108
rect 275060 326068 275066 326080
rect 275830 326068 275836 326080
rect 275888 326068 275894 326120
rect 284754 326068 284760 326120
rect 284812 326108 284818 326120
rect 285030 326108 285036 326120
rect 284812 326080 285036 326108
rect 284812 326068 284818 326080
rect 285030 326068 285036 326080
rect 285088 326068 285094 326120
rect 285674 326068 285680 326120
rect 285732 326108 285738 326120
rect 285950 326108 285956 326120
rect 285732 326080 285956 326108
rect 285732 326068 285738 326080
rect 285950 326068 285956 326080
rect 286008 326068 286014 326120
rect 256418 325972 256424 325984
rect 256344 325944 256424 325972
rect 256418 325932 256424 325944
rect 256476 325932 256482 325984
rect 273346 325864 273352 325916
rect 273404 325904 273410 325916
rect 273898 325904 273904 325916
rect 273404 325876 273904 325904
rect 273404 325864 273410 325876
rect 273898 325864 273904 325876
rect 273956 325864 273962 325916
rect 279050 325796 279056 325848
rect 279108 325836 279114 325848
rect 279326 325836 279332 325848
rect 279108 325808 279332 325836
rect 279108 325796 279114 325808
rect 279326 325796 279332 325808
rect 279384 325796 279390 325848
rect 279510 325728 279516 325780
rect 279568 325728 279574 325780
rect 278774 325524 278780 325576
rect 278832 325564 278838 325576
rect 279418 325564 279424 325576
rect 278832 325536 279424 325564
rect 278832 325524 278838 325536
rect 279418 325524 279424 325536
rect 279476 325524 279482 325576
rect 278774 325388 278780 325440
rect 278832 325428 278838 325440
rect 279528 325428 279556 325728
rect 278832 325400 279556 325428
rect 278832 325388 278838 325400
rect 275646 324980 275652 325032
rect 275704 325020 275710 325032
rect 376754 325020 376760 325032
rect 275704 324992 376760 325020
rect 275704 324980 275710 324992
rect 376754 324980 376760 324992
rect 376812 324980 376818 325032
rect 280890 324912 280896 324964
rect 280948 324952 280954 324964
rect 456794 324952 456800 324964
rect 280948 324924 456800 324952
rect 280948 324912 280954 324924
rect 456794 324912 456800 324924
rect 456852 324912 456858 324964
rect 259730 324164 259736 324216
rect 259788 324204 259794 324216
rect 260558 324204 260564 324216
rect 259788 324176 260564 324204
rect 259788 324164 259794 324176
rect 260558 324164 260564 324176
rect 260616 324164 260622 324216
rect 14 323552 20 323604
rect 72 323592 78 323604
rect 244826 323592 244832 323604
rect 72 323564 244832 323592
rect 72 323552 78 323564
rect 244826 323552 244832 323564
rect 244884 323552 244890 323604
rect 276934 323552 276940 323604
rect 276992 323592 276998 323604
rect 396074 323592 396080 323604
rect 276992 323564 396080 323592
rect 276992 323552 276998 323564
rect 396074 323552 396080 323564
rect 396132 323552 396138 323604
rect 258534 323008 258540 323060
rect 258592 323048 258598 323060
rect 258718 323048 258724 323060
rect 258592 323020 258724 323048
rect 258592 323008 258598 323020
rect 258718 323008 258724 323020
rect 258776 323008 258782 323060
rect 261018 323008 261024 323060
rect 261076 323048 261082 323060
rect 262122 323048 262128 323060
rect 261076 323020 262128 323048
rect 261076 323008 261082 323020
rect 262122 323008 262128 323020
rect 262180 323008 262186 323060
rect 281810 322600 281816 322652
rect 281868 322640 281874 322652
rect 282546 322640 282552 322652
rect 281868 322612 282552 322640
rect 281868 322600 281874 322612
rect 282546 322600 282552 322612
rect 282604 322600 282610 322652
rect 191834 320832 191840 320884
rect 191892 320872 191898 320884
rect 260190 320872 260196 320884
rect 191892 320844 260196 320872
rect 191892 320832 191898 320844
rect 260190 320832 260196 320844
rect 260248 320832 260254 320884
rect 523678 320832 523684 320884
rect 523736 320872 523742 320884
rect 580258 320872 580264 320884
rect 523736 320844 580264 320872
rect 523736 320832 523742 320844
rect 580258 320832 580264 320844
rect 580316 320832 580322 320884
rect 247126 320764 247132 320816
rect 247184 320804 247190 320816
rect 247310 320804 247316 320816
rect 247184 320776 247316 320804
rect 247184 320764 247190 320776
rect 247310 320764 247316 320776
rect 247368 320764 247374 320816
rect 235442 320192 235448 320204
rect 234632 320164 235448 320192
rect 3142 320084 3148 320136
rect 3200 320124 3206 320136
rect 234632 320124 234660 320164
rect 235442 320152 235448 320164
rect 235500 320192 235506 320204
rect 245102 320192 245108 320204
rect 235500 320164 245108 320192
rect 235500 320152 235506 320164
rect 245102 320152 245108 320164
rect 245160 320152 245166 320204
rect 3200 320096 234660 320124
rect 3200 320084 3206 320096
rect 578142 313216 578148 313268
rect 578200 313256 578206 313268
rect 580074 313256 580080 313268
rect 578200 313228 580080 313256
rect 578200 313216 578206 313228
rect 580074 313216 580080 313228
rect 580132 313216 580138 313268
rect 3326 306280 3332 306332
rect 3384 306320 3390 306332
rect 233786 306320 233792 306332
rect 3384 306292 233792 306320
rect 3384 306280 3390 306292
rect 233786 306280 233792 306292
rect 233844 306280 233850 306332
rect 301866 302880 301872 302932
rect 301924 302920 301930 302932
rect 345106 302920 345112 302932
rect 301924 302892 345112 302920
rect 301924 302880 301930 302892
rect 345106 302880 345112 302892
rect 345164 302880 345170 302932
rect 3234 293904 3240 293956
rect 3292 293944 3298 293956
rect 235350 293944 235356 293956
rect 3292 293916 235356 293944
rect 3292 293904 3298 293916
rect 235350 293904 235356 293916
rect 235408 293904 235414 293956
rect 578050 273164 578056 273216
rect 578108 273204 578114 273216
rect 580074 273204 580080 273216
rect 578108 273176 580080 273204
rect 578108 273164 578114 273176
rect 580074 273164 580080 273176
rect 580132 273164 580138 273216
rect 3326 266976 3332 267028
rect 3384 267016 3390 267028
rect 232498 267016 232504 267028
rect 3384 266988 232504 267016
rect 3384 266976 3390 266988
rect 232498 266976 232504 266988
rect 232556 266976 232562 267028
rect 300486 262828 300492 262880
rect 300544 262868 300550 262880
rect 345198 262868 345204 262880
rect 300544 262840 345204 262868
rect 300544 262828 300550 262840
rect 345198 262828 345204 262840
rect 345256 262828 345262 262880
rect 290734 260108 290740 260160
rect 290792 260148 290798 260160
rect 442994 260148 443000 260160
rect 290792 260120 443000 260148
rect 290792 260108 290798 260120
rect 442994 260108 443000 260120
rect 443052 260108 443058 260160
rect 577958 259360 577964 259412
rect 578016 259400 578022 259412
rect 580074 259400 580080 259412
rect 578016 259372 580080 259400
rect 578016 259360 578022 259372
rect 580074 259360 580080 259372
rect 580132 259360 580138 259412
rect 3326 255212 3332 255264
rect 3384 255252 3390 255264
rect 91738 255252 91744 255264
rect 3384 255224 91744 255252
rect 3384 255212 3390 255224
rect 91738 255212 91744 255224
rect 91796 255212 91802 255264
rect 3326 241408 3332 241460
rect 3384 241448 3390 241460
rect 90450 241448 90456 241460
rect 3384 241420 90456 241448
rect 3384 241408 3390 241420
rect 90450 241408 90456 241420
rect 90508 241408 90514 241460
rect 577774 219172 577780 219224
rect 577832 219212 577838 219224
rect 579706 219212 579712 219224
rect 577832 219184 579712 219212
rect 577832 219172 577838 219184
rect 579706 219172 579712 219184
rect 579764 219172 579770 219224
rect 3326 214548 3332 214600
rect 3384 214588 3390 214600
rect 237466 214588 237472 214600
rect 3384 214560 237472 214588
rect 3384 214548 3390 214560
rect 237466 214548 237472 214560
rect 237524 214548 237530 214600
rect 287606 193808 287612 193860
rect 287664 193848 287670 193860
rect 547874 193848 547880 193860
rect 287664 193820 547880 193848
rect 287664 193808 287670 193820
rect 547874 193808 547880 193820
rect 547932 193808 547938 193860
rect 154574 191088 154580 191140
rect 154632 191128 154638 191140
rect 257062 191128 257068 191140
rect 154632 191100 257068 191128
rect 154632 191088 154638 191100
rect 257062 191088 257068 191100
rect 257120 191088 257126 191140
rect 294598 184220 294604 184272
rect 294656 184260 294662 184272
rect 449894 184260 449900 184272
rect 294656 184232 449900 184260
rect 294656 184220 294662 184232
rect 449894 184220 449900 184232
rect 449952 184220 449958 184272
rect 282178 184152 282184 184204
rect 282236 184192 282242 184204
rect 471974 184192 471980 184204
rect 282236 184164 471980 184192
rect 282236 184152 282242 184164
rect 471974 184152 471980 184164
rect 472032 184152 472038 184204
rect 277946 180140 277952 180192
rect 278004 180180 278010 180192
rect 418154 180180 418160 180192
rect 278004 180152 418160 180180
rect 278004 180140 278010 180152
rect 418154 180140 418160 180152
rect 418212 180140 418218 180192
rect 290182 180072 290188 180124
rect 290240 180112 290246 180124
rect 580994 180112 581000 180124
rect 290240 180084 581000 180112
rect 290240 180072 290246 180084
rect 580994 180072 581000 180084
rect 581052 180072 581058 180124
rect 577866 179324 577872 179376
rect 577924 179364 577930 179376
rect 579706 179364 579712 179376
rect 577924 179336 579712 179364
rect 577924 179324 577930 179336
rect 579706 179324 579712 179336
rect 579764 179324 579770 179376
rect 160186 179120 160192 179172
rect 160244 179160 160250 179172
rect 256970 179160 256976 179172
rect 160244 179132 256976 179160
rect 160244 179120 160250 179132
rect 256970 179120 256976 179132
rect 257028 179120 257034 179172
rect 115934 179052 115940 179104
rect 115992 179092 115998 179104
rect 254394 179092 254400 179104
rect 115992 179064 254400 179092
rect 115992 179052 115998 179064
rect 254394 179052 254400 179064
rect 254452 179052 254458 179104
rect 273806 179052 273812 179104
rect 273864 179092 273870 179104
rect 368474 179092 368480 179104
rect 273864 179064 368480 179092
rect 273864 179052 273870 179064
rect 368474 179052 368480 179064
rect 368532 179052 368538 179104
rect 109034 178984 109040 179036
rect 109092 179024 109098 179036
rect 253290 179024 253296 179036
rect 109092 178996 253296 179024
rect 109092 178984 109098 178996
rect 253290 178984 253296 178996
rect 253348 178984 253354 179036
rect 283558 178984 283564 179036
rect 283616 179024 283622 179036
rect 386414 179024 386420 179036
rect 283616 178996 386420 179024
rect 283616 178984 283622 178996
rect 386414 178984 386420 178996
rect 386472 178984 386478 179036
rect 104894 178916 104900 178968
rect 104952 178956 104958 178968
rect 253198 178956 253204 178968
rect 104952 178928 253204 178956
rect 104952 178916 104958 178928
rect 253198 178916 253204 178928
rect 253256 178916 253262 178968
rect 277854 178916 277860 178968
rect 277912 178956 277918 178968
rect 415394 178956 415400 178968
rect 277912 178928 415400 178956
rect 277912 178916 277918 178928
rect 415394 178916 415400 178928
rect 415452 178916 415458 178968
rect 97994 178848 98000 178900
rect 98052 178888 98058 178900
rect 253106 178888 253112 178900
rect 98052 178860 253112 178888
rect 98052 178848 98058 178860
rect 253106 178848 253112 178860
rect 253164 178848 253170 178900
rect 288894 178848 288900 178900
rect 288952 178888 288958 178900
rect 560294 178888 560300 178900
rect 288952 178860 560300 178888
rect 288952 178848 288958 178860
rect 560294 178848 560300 178860
rect 560352 178848 560358 178900
rect 67634 178780 67640 178832
rect 67692 178820 67698 178832
rect 250530 178820 250536 178832
rect 67692 178792 250536 178820
rect 67692 178780 67698 178792
rect 250530 178780 250536 178792
rect 250588 178780 250594 178832
rect 288802 178780 288808 178832
rect 288860 178820 288866 178832
rect 567194 178820 567200 178832
rect 288860 178792 567200 178820
rect 288860 178780 288866 178792
rect 567194 178780 567200 178792
rect 567252 178780 567258 178832
rect 49694 178712 49700 178764
rect 49752 178752 49758 178764
rect 248874 178752 248880 178764
rect 49752 178724 248880 178752
rect 49752 178712 49758 178724
rect 248874 178712 248880 178724
rect 248932 178712 248938 178764
rect 289998 178712 290004 178764
rect 290056 178752 290062 178764
rect 574094 178752 574100 178764
rect 290056 178724 574100 178752
rect 290056 178712 290062 178724
rect 574094 178712 574100 178724
rect 574152 178712 574158 178764
rect 2774 178644 2780 178696
rect 2832 178684 2838 178696
rect 244458 178684 244464 178696
rect 2832 178656 244464 178684
rect 2832 178644 2838 178656
rect 244458 178644 244464 178656
rect 244516 178644 244522 178696
rect 290090 178644 290096 178696
rect 290148 178684 290154 178696
rect 578234 178684 578240 178696
rect 290148 178656 578240 178684
rect 290148 178644 290154 178656
rect 578234 178644 578240 178656
rect 578292 178644 578298 178696
rect 176654 177828 176660 177880
rect 176712 177868 176718 177880
rect 258442 177868 258448 177880
rect 176712 177840 258448 177868
rect 176712 177828 176718 177840
rect 258442 177828 258448 177840
rect 258500 177828 258506 177880
rect 162854 177760 162860 177812
rect 162912 177800 162918 177812
rect 257154 177800 257160 177812
rect 162912 177772 257160 177800
rect 162912 177760 162918 177772
rect 257154 177760 257160 177772
rect 257212 177760 257218 177812
rect 280706 177760 280712 177812
rect 280764 177800 280770 177812
rect 452654 177800 452660 177812
rect 280764 177772 452660 177800
rect 280764 177760 280770 177772
rect 452654 177760 452660 177772
rect 452712 177760 452718 177812
rect 158714 177692 158720 177744
rect 158772 177732 158778 177744
rect 256878 177732 256884 177744
rect 158772 177704 256884 177732
rect 158772 177692 158778 177704
rect 256878 177692 256884 177704
rect 256936 177692 256942 177744
rect 280798 177692 280804 177744
rect 280856 177732 280862 177744
rect 459554 177732 459560 177744
rect 280856 177704 459560 177732
rect 280856 177692 280862 177704
rect 459554 177692 459560 177704
rect 459612 177692 459618 177744
rect 151906 177624 151912 177676
rect 151964 177664 151970 177676
rect 257430 177664 257436 177676
rect 151964 177636 257436 177664
rect 151964 177624 151970 177636
rect 257430 177624 257436 177636
rect 257488 177624 257494 177676
rect 284846 177624 284852 177676
rect 284904 177664 284910 177676
rect 503714 177664 503720 177676
rect 284904 177636 503720 177664
rect 284904 177624 284910 177636
rect 503714 177624 503720 177636
rect 503772 177624 503778 177676
rect 144914 177556 144920 177608
rect 144972 177596 144978 177608
rect 255682 177596 255688 177608
rect 144972 177568 255688 177596
rect 144972 177556 144978 177568
rect 255682 177556 255688 177568
rect 255740 177556 255746 177608
rect 284938 177556 284944 177608
rect 284996 177596 285002 177608
rect 510614 177596 510620 177608
rect 284996 177568 510620 177596
rect 284996 177556 285002 177568
rect 510614 177556 510620 177568
rect 510672 177556 510678 177608
rect 66254 177488 66260 177540
rect 66312 177528 66318 177540
rect 250438 177528 250444 177540
rect 66312 177500 250444 177528
rect 66312 177488 66318 177500
rect 250438 177488 250444 177500
rect 250496 177488 250502 177540
rect 286134 177488 286140 177540
rect 286192 177528 286198 177540
rect 521654 177528 521660 177540
rect 286192 177500 521660 177528
rect 286192 177488 286198 177500
rect 521654 177488 521660 177500
rect 521712 177488 521718 177540
rect 55214 177420 55220 177472
rect 55272 177460 55278 177472
rect 248782 177460 248788 177472
rect 55272 177432 248788 177460
rect 55272 177420 55278 177432
rect 248782 177420 248788 177432
rect 248840 177420 248846 177472
rect 286042 177420 286048 177472
rect 286100 177460 286106 177472
rect 524414 177460 524420 177472
rect 286100 177432 524420 177460
rect 286100 177420 286106 177432
rect 524414 177420 524420 177432
rect 524472 177420 524478 177472
rect 48314 177352 48320 177404
rect 48372 177392 48378 177404
rect 248690 177392 248696 177404
rect 48372 177364 248696 177392
rect 48372 177352 48378 177364
rect 248690 177352 248696 177364
rect 248748 177352 248754 177404
rect 287514 177352 287520 177404
rect 287572 177392 287578 177404
rect 542354 177392 542360 177404
rect 287572 177364 542360 177392
rect 287572 177352 287578 177364
rect 542354 177352 542360 177364
rect 542412 177352 542418 177404
rect 17954 177284 17960 177336
rect 18012 177324 18018 177336
rect 246114 177324 246120 177336
rect 18012 177296 246120 177324
rect 18012 177284 18018 177296
rect 246114 177284 246120 177296
rect 246172 177284 246178 177336
rect 287422 177284 287428 177336
rect 287480 177324 287486 177336
rect 546494 177324 546500 177336
rect 287480 177296 546500 177324
rect 287480 177284 287486 177296
rect 546494 177284 546500 177296
rect 546552 177284 546558 177336
rect 275370 176400 275376 176452
rect 275428 176440 275434 176452
rect 382274 176440 382280 176452
rect 275428 176412 382280 176440
rect 275428 176400 275434 176412
rect 382274 176400 382280 176412
rect 382332 176400 382338 176452
rect 275186 176332 275192 176384
rect 275244 176372 275250 176384
rect 385034 176372 385040 176384
rect 275244 176344 385040 176372
rect 275244 176332 275250 176344
rect 385034 176332 385040 176344
rect 385092 176332 385098 176384
rect 275278 176264 275284 176316
rect 275336 176304 275342 176316
rect 389174 176304 389180 176316
rect 275336 176276 389180 176304
rect 275336 176264 275342 176276
rect 389174 176264 389180 176276
rect 389232 176264 389238 176316
rect 276290 176196 276296 176248
rect 276348 176236 276354 176248
rect 402974 176236 402980 176248
rect 276348 176208 402980 176236
rect 276348 176196 276354 176208
rect 402974 176196 402980 176208
rect 403032 176196 403038 176248
rect 277670 176128 277676 176180
rect 277728 176168 277734 176180
rect 416774 176168 416780 176180
rect 277728 176140 416780 176168
rect 277728 176128 277734 176140
rect 416774 176128 416780 176140
rect 416832 176128 416838 176180
rect 293494 176060 293500 176112
rect 293552 176100 293558 176112
rect 436094 176100 436100 176112
rect 293552 176072 436100 176100
rect 293552 176060 293558 176072
rect 436094 176060 436100 176072
rect 436152 176060 436158 176112
rect 277762 175992 277768 176044
rect 277820 176032 277826 176044
rect 423766 176032 423772 176044
rect 277820 176004 423772 176032
rect 277820 175992 277826 176004
rect 423766 175992 423772 176004
rect 423824 175992 423830 176044
rect 279418 175924 279424 175976
rect 279476 175964 279482 175976
rect 431954 175964 431960 175976
rect 279476 175936 431960 175964
rect 279476 175924 279482 175936
rect 431954 175924 431960 175936
rect 432012 175924 432018 175976
rect 273622 174768 273628 174820
rect 273680 174808 273686 174820
rect 367094 174808 367100 174820
rect 273680 174780 367100 174808
rect 273680 174768 273686 174780
rect 367094 174768 367100 174780
rect 367152 174768 367158 174820
rect 273714 174700 273720 174752
rect 273772 174740 273778 174752
rect 371234 174740 371240 174752
rect 273772 174712 371240 174740
rect 273772 174700 273778 174712
rect 371234 174700 371240 174712
rect 371292 174700 371298 174752
rect 275094 174632 275100 174684
rect 275152 174672 275158 174684
rect 378134 174672 378140 174684
rect 275152 174644 378140 174672
rect 275152 174632 275158 174644
rect 378134 174632 378140 174644
rect 378192 174632 378198 174684
rect 280614 174564 280620 174616
rect 280672 174604 280678 174616
rect 454034 174604 454040 174616
rect 280672 174576 454040 174604
rect 280672 174564 280678 174576
rect 454034 174564 454040 174576
rect 454092 174564 454098 174616
rect 287330 174496 287336 174548
rect 287388 174536 287394 174548
rect 539686 174536 539692 174548
rect 287388 174508 539692 174536
rect 287388 174496 287394 174508
rect 539686 174496 539692 174508
rect 539744 174496 539750 174548
rect 292114 173476 292120 173528
rect 292172 173516 292178 173528
rect 404354 173516 404360 173528
rect 292172 173488 404360 173516
rect 292172 173476 292178 173488
rect 404354 173476 404360 173488
rect 404412 173476 404418 173528
rect 285858 173408 285864 173460
rect 285916 173448 285922 173460
rect 520274 173448 520280 173460
rect 285916 173420 520280 173448
rect 285916 173408 285922 173420
rect 520274 173408 520280 173420
rect 520332 173408 520338 173460
rect 285950 173340 285956 173392
rect 286008 173380 286014 173392
rect 527174 173380 527180 173392
rect 286008 173352 527180 173380
rect 286008 173340 286014 173352
rect 527174 173340 527180 173352
rect 527232 173340 527238 173392
rect 287238 173272 287244 173324
rect 287296 173312 287302 173324
rect 540974 173312 540980 173324
rect 287296 173284 540980 173312
rect 287296 173272 287302 173284
rect 540974 173272 540980 173284
rect 541032 173272 541038 173324
rect 288710 173204 288716 173256
rect 288768 173244 288774 173256
rect 563054 173244 563060 173256
rect 288768 173216 563060 173244
rect 288768 173204 288774 173216
rect 563054 173204 563060 173216
rect 563112 173204 563118 173256
rect 289906 173136 289912 173188
rect 289964 173176 289970 173188
rect 576854 173176 576860 173188
rect 289964 173148 576860 173176
rect 289964 173136 289970 173148
rect 576854 173136 576860 173148
rect 576912 173136 576918 173188
rect 291930 172320 291936 172372
rect 291988 172360 291994 172372
rect 393314 172360 393320 172372
rect 291988 172332 393320 172360
rect 291988 172320 291994 172332
rect 393314 172320 393320 172332
rect 393372 172320 393378 172372
rect 292022 172252 292028 172304
rect 292080 172292 292086 172304
rect 397454 172292 397460 172304
rect 292080 172264 397460 172292
rect 292080 172252 292086 172264
rect 397454 172252 397460 172264
rect 397512 172252 397518 172304
rect 295978 172184 295984 172236
rect 296036 172224 296042 172236
rect 456886 172224 456892 172236
rect 296036 172196 456892 172224
rect 296036 172184 296042 172196
rect 456886 172184 456892 172196
rect 456944 172184 456950 172236
rect 283466 172116 283472 172168
rect 283524 172156 283530 172168
rect 484394 172156 484400 172168
rect 283524 172128 484400 172156
rect 283524 172116 283530 172128
rect 484394 172116 484400 172128
rect 484452 172116 484458 172168
rect 283282 172048 283288 172100
rect 283340 172088 283346 172100
rect 488534 172088 488540 172100
rect 283340 172060 488540 172088
rect 283340 172048 283346 172060
rect 488534 172048 488540 172060
rect 488592 172048 488598 172100
rect 283190 171980 283196 172032
rect 283248 172020 283254 172032
rect 490006 172020 490012 172032
rect 283248 171992 490012 172020
rect 283248 171980 283254 171992
rect 490006 171980 490012 171992
rect 490064 171980 490070 172032
rect 283374 171912 283380 171964
rect 283432 171952 283438 171964
rect 492674 171952 492680 171964
rect 283432 171924 492680 171952
rect 283432 171912 283438 171924
rect 492674 171912 492680 171924
rect 492732 171912 492738 171964
rect 284662 171844 284668 171896
rect 284720 171884 284726 171896
rect 506474 171884 506480 171896
rect 284720 171856 506480 171884
rect 284720 171844 284726 171856
rect 506474 171844 506480 171856
rect 506532 171844 506538 171896
rect 284754 171776 284760 171828
rect 284812 171816 284818 171828
rect 513374 171816 513380 171828
rect 284812 171788 513380 171816
rect 284812 171776 284818 171788
rect 513374 171776 513380 171788
rect 513432 171776 513438 171828
rect 276750 170756 276756 170808
rect 276808 170796 276814 170808
rect 364334 170796 364340 170808
rect 276808 170768 364340 170796
rect 276808 170756 276814 170768
rect 364334 170756 364340 170768
rect 364392 170756 364398 170808
rect 293402 170688 293408 170740
rect 293460 170728 293466 170740
rect 422294 170728 422300 170740
rect 293460 170700 422300 170728
rect 293460 170688 293466 170700
rect 422294 170688 422300 170700
rect 422352 170688 422358 170740
rect 279142 170620 279148 170672
rect 279200 170660 279206 170672
rect 432046 170660 432052 170672
rect 279200 170632 432052 170660
rect 279200 170620 279206 170632
rect 432046 170620 432052 170632
rect 432104 170620 432110 170672
rect 279234 170552 279240 170604
rect 279292 170592 279298 170604
rect 434714 170592 434720 170604
rect 279292 170564 434720 170592
rect 279292 170552 279298 170564
rect 434714 170552 434720 170564
rect 434772 170552 434778 170604
rect 279326 170484 279332 170536
rect 279384 170524 279390 170536
rect 441614 170524 441620 170536
rect 279384 170496 441620 170524
rect 279384 170484 279390 170496
rect 441614 170484 441620 170496
rect 441672 170484 441678 170536
rect 281994 170416 282000 170468
rect 282052 170456 282058 170468
rect 473354 170456 473360 170468
rect 282052 170428 473360 170456
rect 282052 170416 282058 170428
rect 473354 170416 473360 170428
rect 473412 170416 473418 170468
rect 282086 170348 282092 170400
rect 282144 170388 282150 170400
rect 476114 170388 476120 170400
rect 282144 170360 476120 170388
rect 282144 170348 282150 170360
rect 476114 170348 476120 170360
rect 476172 170348 476178 170400
rect 273898 169192 273904 169244
rect 273956 169232 273962 169244
rect 349338 169232 349344 169244
rect 273956 169204 349344 169232
rect 273956 169192 273962 169204
rect 349338 169192 349344 169204
rect 349396 169192 349402 169244
rect 280522 169124 280528 169176
rect 280580 169164 280586 169176
rect 462314 169164 462320 169176
rect 280580 169136 462320 169164
rect 280580 169124 280586 169136
rect 462314 169124 462320 169136
rect 462372 169124 462378 169176
rect 281902 169056 281908 169108
rect 281960 169096 281966 169108
rect 469214 169096 469220 169108
rect 281960 169068 469220 169096
rect 281960 169056 281966 169068
rect 469214 169056 469220 169068
rect 469272 169056 469278 169108
rect 283098 168988 283104 169040
rect 283156 169028 283162 169040
rect 485774 169028 485780 169040
rect 283156 169000 485780 169028
rect 283156 168988 283162 169000
rect 485774 168988 485780 169000
rect 485832 168988 485838 169040
rect 278866 168104 278872 168156
rect 278924 168144 278930 168156
rect 433334 168144 433340 168156
rect 278924 168116 433340 168144
rect 278924 168104 278930 168116
rect 433334 168104 433340 168116
rect 433392 168104 433398 168156
rect 279050 168036 279056 168088
rect 279108 168076 279114 168088
rect 437474 168076 437480 168088
rect 279108 168048 437480 168076
rect 279108 168036 279114 168048
rect 437474 168036 437480 168048
rect 437532 168036 437538 168088
rect 278958 167968 278964 168020
rect 279016 168008 279022 168020
rect 440234 168008 440240 168020
rect 279016 167980 440240 168008
rect 279016 167968 279022 167980
rect 440234 167968 440240 167980
rect 440292 167968 440298 168020
rect 280338 167900 280344 167952
rect 280396 167940 280402 167952
rect 455414 167940 455420 167952
rect 280396 167912 455420 167940
rect 280396 167900 280402 167912
rect 455414 167900 455420 167912
rect 455472 167900 455478 167952
rect 280430 167832 280436 167884
rect 280488 167872 280494 167884
rect 458174 167872 458180 167884
rect 280488 167844 458180 167872
rect 280488 167832 280494 167844
rect 458174 167832 458180 167844
rect 458232 167832 458238 167884
rect 280246 167764 280252 167816
rect 280304 167804 280310 167816
rect 460934 167804 460940 167816
rect 280304 167776 460940 167804
rect 280304 167764 280310 167776
rect 460934 167764 460940 167776
rect 460992 167764 460998 167816
rect 281810 167696 281816 167748
rect 281868 167736 281874 167748
rect 478874 167736 478880 167748
rect 281868 167708 478880 167736
rect 281868 167696 281874 167708
rect 478874 167696 478880 167708
rect 478932 167696 478938 167748
rect 289814 167628 289820 167680
rect 289872 167668 289878 167680
rect 582374 167668 582380 167680
rect 289872 167640 582380 167668
rect 289872 167628 289878 167640
rect 582374 167628 582380 167640
rect 582432 167628 582438 167680
rect 407758 166948 407764 167000
rect 407816 166988 407822 167000
rect 580166 166988 580172 167000
rect 407816 166960 580172 166988
rect 407816 166948 407822 166960
rect 580166 166948 580172 166960
rect 580224 166948 580230 167000
rect 277578 166608 277584 166660
rect 277636 166648 277642 166660
rect 412634 166648 412640 166660
rect 277636 166620 412640 166648
rect 277636 166608 277642 166620
rect 412634 166608 412640 166620
rect 412692 166608 412698 166660
rect 293310 166540 293316 166592
rect 293368 166580 293374 166592
rect 429194 166580 429200 166592
rect 293368 166552 429200 166580
rect 293368 166540 293374 166552
rect 429194 166540 429200 166552
rect 429252 166540 429258 166592
rect 277394 166472 277400 166524
rect 277452 166512 277458 166524
rect 415486 166512 415492 166524
rect 277452 166484 415492 166512
rect 277452 166472 277458 166484
rect 415486 166472 415492 166484
rect 415544 166472 415550 166524
rect 277486 166404 277492 166456
rect 277544 166444 277550 166456
rect 419534 166444 419540 166456
rect 277544 166416 419540 166444
rect 277544 166404 277550 166416
rect 419534 166404 419540 166416
rect 419592 166404 419598 166456
rect 278774 166336 278780 166388
rect 278832 166376 278838 166388
rect 440326 166376 440332 166388
rect 278832 166348 440332 166376
rect 278832 166336 278838 166348
rect 440326 166336 440332 166348
rect 440384 166336 440390 166388
rect 291838 166268 291844 166320
rect 291896 166308 291902 166320
rect 554774 166308 554780 166320
rect 291896 166280 554780 166308
rect 291896 166268 291902 166280
rect 554774 166268 554780 166280
rect 554832 166268 554838 166320
rect 274726 165248 274732 165300
rect 274784 165288 274790 165300
rect 382366 165288 382372 165300
rect 274784 165260 382372 165288
rect 274784 165248 274790 165260
rect 382366 165248 382372 165260
rect 382424 165248 382430 165300
rect 274818 165180 274824 165232
rect 274876 165220 274882 165232
rect 383654 165220 383660 165232
rect 274876 165192 383660 165220
rect 274876 165180 274882 165192
rect 383654 165180 383660 165192
rect 383712 165180 383718 165232
rect 274910 165112 274916 165164
rect 274968 165152 274974 165164
rect 387794 165152 387800 165164
rect 274968 165124 387800 165152
rect 274968 165112 274974 165124
rect 387794 165112 387800 165124
rect 387852 165112 387858 165164
rect 275002 165044 275008 165096
rect 275060 165084 275066 165096
rect 390646 165084 390652 165096
rect 275060 165056 390652 165084
rect 275060 165044 275066 165056
rect 390646 165044 390652 165056
rect 390704 165044 390710 165096
rect 276198 164976 276204 165028
rect 276256 165016 276262 165028
rect 400214 165016 400220 165028
rect 276256 164988 400220 165016
rect 276256 164976 276262 164988
rect 400214 164976 400220 164988
rect 400272 164976 400278 165028
rect 276106 164908 276112 164960
rect 276164 164948 276170 164960
rect 401594 164948 401600 164960
rect 276164 164920 401600 164948
rect 276164 164908 276170 164920
rect 401594 164908 401600 164920
rect 401652 164908 401658 164960
rect 276014 164840 276020 164892
rect 276072 164880 276078 164892
rect 405734 164880 405740 164892
rect 276072 164852 405740 164880
rect 276072 164840 276078 164852
rect 405734 164840 405740 164852
rect 405792 164840 405798 164892
rect 3326 164160 3332 164212
rect 3384 164200 3390 164212
rect 234798 164200 234804 164212
rect 3384 164172 234804 164200
rect 3384 164160 3390 164172
rect 234798 164160 234804 164172
rect 234856 164160 234862 164212
rect 273438 163888 273444 163940
rect 273496 163928 273502 163940
rect 362954 163928 362960 163940
rect 273496 163900 362960 163928
rect 273496 163888 273502 163900
rect 362954 163888 362960 163900
rect 363012 163888 363018 163940
rect 273346 163820 273352 163872
rect 273404 163860 273410 163872
rect 365806 163860 365812 163872
rect 273404 163832 365812 163860
rect 273404 163820 273410 163832
rect 365806 163820 365812 163832
rect 365864 163820 365870 163872
rect 273530 163752 273536 163804
rect 273588 163792 273594 163804
rect 369854 163792 369860 163804
rect 273588 163764 369860 163792
rect 273588 163752 273594 163764
rect 369854 163752 369860 163764
rect 369912 163752 369918 163804
rect 256418 163684 256424 163736
rect 256476 163724 256482 163736
rect 357434 163724 357440 163736
rect 256476 163696 357440 163724
rect 256476 163684 256482 163696
rect 357434 163684 357440 163696
rect 357492 163684 357498 163736
rect 274634 163616 274640 163668
rect 274692 163656 274698 163668
rect 380894 163656 380900 163668
rect 274692 163628 380900 163656
rect 274692 163616 274698 163628
rect 380894 163616 380900 163628
rect 380952 163616 380958 163668
rect 311158 163548 311164 163600
rect 311216 163588 311222 163600
rect 581086 163588 581092 163600
rect 311216 163560 581092 163588
rect 311216 163548 311222 163560
rect 581086 163548 581092 163560
rect 581144 163548 581150 163600
rect 234798 163480 234804 163532
rect 234856 163520 234862 163532
rect 235534 163520 235540 163532
rect 234856 163492 235540 163520
rect 234856 163480 234862 163492
rect 235534 163480 235540 163492
rect 235592 163520 235598 163532
rect 272610 163520 272616 163532
rect 235592 163492 272616 163520
rect 235592 163480 235598 163492
rect 272610 163480 272616 163492
rect 272668 163480 272674 163532
rect 288618 163480 288624 163532
rect 288676 163520 288682 163532
rect 558914 163520 558920 163532
rect 288676 163492 558920 163520
rect 288676 163480 288682 163492
rect 558914 163480 558920 163492
rect 558972 163480 558978 163532
rect 276658 162256 276664 162308
rect 276716 162296 276722 162308
rect 372614 162296 372620 162308
rect 276716 162268 372620 162296
rect 276716 162256 276722 162268
rect 372614 162256 372620 162268
rect 372672 162256 372678 162308
rect 284570 162188 284576 162240
rect 284628 162228 284634 162240
rect 506566 162228 506572 162240
rect 284628 162200 506572 162228
rect 284628 162188 284634 162200
rect 506566 162188 506572 162200
rect 506624 162188 506630 162240
rect 272610 162120 272616 162172
rect 272668 162160 272674 162172
rect 285766 162160 285772 162172
rect 272668 162132 285772 162160
rect 272668 162120 272674 162132
rect 285766 162120 285772 162132
rect 285824 162120 285830 162172
rect 288526 162120 288532 162172
rect 288584 162160 288590 162172
rect 564526 162160 564532 162172
rect 288584 162132 564532 162160
rect 288584 162120 288590 162132
rect 564526 162120 564532 162132
rect 564584 162120 564590 162172
rect 242618 161372 242624 161424
rect 242676 161412 242682 161424
rect 266998 161412 267004 161424
rect 242676 161384 267004 161412
rect 242676 161372 242682 161384
rect 266998 161372 267004 161384
rect 267056 161372 267062 161424
rect 245470 161304 245476 161356
rect 245528 161344 245534 161356
rect 269942 161344 269948 161356
rect 245528 161316 269948 161344
rect 245528 161304 245534 161316
rect 269942 161304 269948 161316
rect 270000 161304 270006 161356
rect 259546 161236 259552 161288
rect 259604 161276 259610 161288
rect 299474 161276 299480 161288
rect 259604 161248 299480 161276
rect 259604 161236 259610 161248
rect 299474 161236 299480 161248
rect 299532 161236 299538 161288
rect 242710 161168 242716 161220
rect 242768 161208 242774 161220
rect 267182 161208 267188 161220
rect 242768 161180 267188 161208
rect 242768 161168 242774 161180
rect 267182 161168 267188 161180
rect 267240 161168 267246 161220
rect 272518 161168 272524 161220
rect 272576 161208 272582 161220
rect 347958 161208 347964 161220
rect 272576 161180 347964 161208
rect 272576 161168 272582 161180
rect 347958 161168 347964 161180
rect 348016 161168 348022 161220
rect 243998 161100 244004 161152
rect 244056 161140 244062 161152
rect 268562 161140 268568 161152
rect 244056 161112 268568 161140
rect 244056 161100 244062 161112
rect 268562 161100 268568 161112
rect 268620 161100 268626 161152
rect 271230 161100 271236 161152
rect 271288 161140 271294 161152
rect 348234 161140 348240 161152
rect 271288 161112 348240 161140
rect 271288 161100 271294 161112
rect 348234 161100 348240 161112
rect 348292 161100 348298 161152
rect 242066 161032 242072 161084
rect 242124 161072 242130 161084
rect 267090 161072 267096 161084
rect 242124 161044 267096 161072
rect 242124 161032 242130 161044
rect 267090 161032 267096 161044
rect 267148 161032 267154 161084
rect 272426 161032 272432 161084
rect 272484 161072 272490 161084
rect 350534 161072 350540 161084
rect 272484 161044 350540 161072
rect 272484 161032 272490 161044
rect 350534 161032 350540 161044
rect 350592 161032 350598 161084
rect 241330 160964 241336 161016
rect 241388 161004 241394 161016
rect 268010 161004 268016 161016
rect 241388 160976 268016 161004
rect 241388 160964 241394 160976
rect 268010 160964 268016 160976
rect 268068 160964 268074 161016
rect 281442 160964 281448 161016
rect 281500 161004 281506 161016
rect 448606 161004 448612 161016
rect 281500 160976 448612 161004
rect 281500 160964 281506 160976
rect 448606 160964 448612 160976
rect 448664 160964 448670 161016
rect 239950 160896 239956 160948
rect 240008 160936 240014 160948
rect 268286 160936 268292 160948
rect 240008 160908 268292 160936
rect 240008 160896 240014 160908
rect 268286 160896 268292 160908
rect 268344 160896 268350 160948
rect 281718 160896 281724 160948
rect 281776 160936 281782 160948
rect 477494 160936 477500 160948
rect 281776 160908 477500 160936
rect 281776 160896 281782 160908
rect 477494 160896 477500 160908
rect 477552 160896 477558 160948
rect 239674 160828 239680 160880
rect 239732 160868 239738 160880
rect 268102 160868 268108 160880
rect 239732 160840 268108 160868
rect 239732 160828 239738 160840
rect 268102 160828 268108 160840
rect 268160 160828 268166 160880
rect 287146 160828 287152 160880
rect 287204 160868 287210 160880
rect 543734 160868 543740 160880
rect 287204 160840 543740 160868
rect 287204 160828 287210 160840
rect 543734 160828 543740 160840
rect 543792 160828 543798 160880
rect 239766 160760 239772 160812
rect 239824 160800 239830 160812
rect 268470 160800 268476 160812
rect 239824 160772 268476 160800
rect 239824 160760 239830 160772
rect 268470 160760 268476 160772
rect 268528 160760 268534 160812
rect 287054 160760 287060 160812
rect 287112 160800 287118 160812
rect 547966 160800 547972 160812
rect 287112 160772 547972 160800
rect 287112 160760 287118 160772
rect 547966 160760 547972 160772
rect 548024 160760 548030 160812
rect 44174 160692 44180 160744
rect 44232 160732 44238 160744
rect 247678 160732 247684 160744
rect 44232 160704 247684 160732
rect 44232 160692 44238 160704
rect 247678 160692 247684 160704
rect 247736 160692 247742 160744
rect 250990 160692 250996 160744
rect 251048 160732 251054 160744
rect 268378 160732 268384 160744
rect 251048 160704 268384 160732
rect 251048 160692 251054 160704
rect 268378 160692 268384 160704
rect 268436 160692 268442 160744
rect 288434 160692 288440 160744
rect 288492 160732 288498 160744
rect 561674 160732 561680 160744
rect 288492 160704 561680 160732
rect 288492 160692 288498 160704
rect 561674 160692 561680 160704
rect 561732 160692 561738 160744
rect 242802 160624 242808 160676
rect 242860 160664 242866 160676
rect 265434 160664 265440 160676
rect 242860 160636 265440 160664
rect 242860 160624 242866 160636
rect 265434 160624 265440 160636
rect 265492 160624 265498 160676
rect 246850 160556 246856 160608
rect 246908 160596 246914 160608
rect 268194 160596 268200 160608
rect 246908 160568 268200 160596
rect 246908 160556 246914 160568
rect 268194 160556 268200 160568
rect 268252 160556 268258 160608
rect 248690 160488 248696 160540
rect 248748 160528 248754 160540
rect 264146 160528 264152 160540
rect 248748 160500 264152 160528
rect 248748 160488 248754 160500
rect 264146 160488 264152 160500
rect 264204 160488 264210 160540
rect 251634 159808 251640 159860
rect 251692 159848 251698 159860
rect 263962 159848 263968 159860
rect 251692 159820 263968 159848
rect 251692 159808 251698 159820
rect 263962 159808 263968 159820
rect 264020 159808 264026 159860
rect 247586 159740 247592 159792
rect 247644 159780 247650 159792
rect 264054 159780 264060 159792
rect 247644 159752 264060 159780
rect 247644 159740 247650 159752
rect 264054 159740 264060 159752
rect 264112 159740 264118 159792
rect 244458 159672 244464 159724
rect 244516 159712 244522 159724
rect 263870 159712 263876 159724
rect 244516 159684 263876 159712
rect 244516 159672 244522 159684
rect 263870 159672 263876 159684
rect 263928 159672 263934 159724
rect 230474 159604 230480 159656
rect 230532 159644 230538 159656
rect 262490 159644 262496 159656
rect 230532 159616 262496 159644
rect 230532 159604 230538 159616
rect 262490 159604 262496 159616
rect 262548 159604 262554 159656
rect 223574 159536 223580 159588
rect 223632 159576 223638 159588
rect 262398 159576 262404 159588
rect 223632 159548 262404 159576
rect 223632 159536 223638 159548
rect 262398 159536 262404 159548
rect 262456 159536 262462 159588
rect 300394 159536 300400 159588
rect 300452 159576 300458 159588
rect 327626 159576 327632 159588
rect 300452 159548 327632 159576
rect 300452 159536 300458 159548
rect 327626 159536 327632 159548
rect 327684 159536 327690 159588
rect 382918 159536 382924 159588
rect 382976 159576 382982 159588
rect 465166 159576 465172 159588
rect 382976 159548 465172 159576
rect 382976 159536 382982 159548
rect 465166 159536 465172 159548
rect 465224 159536 465230 159588
rect 222194 159468 222200 159520
rect 222252 159508 222258 159520
rect 262582 159508 262588 159520
rect 222252 159480 262588 159508
rect 222252 159468 222258 159480
rect 262582 159468 262588 159480
rect 262640 159468 262646 159520
rect 281626 159468 281632 159520
rect 281684 159508 281690 159520
rect 470594 159508 470600 159520
rect 281684 159480 470600 159508
rect 281684 159468 281690 159480
rect 470594 159468 470600 159480
rect 470652 159468 470658 159520
rect 212534 159400 212540 159452
rect 212592 159440 212598 159452
rect 261294 159440 261300 159452
rect 212592 159412 261300 159440
rect 212592 159400 212598 159412
rect 261294 159400 261300 159412
rect 261352 159400 261358 159452
rect 286686 159400 286692 159452
rect 286744 159440 286750 159452
rect 525794 159440 525800 159452
rect 286744 159412 525800 159440
rect 286744 159400 286750 159412
rect 525794 159400 525800 159412
rect 525852 159400 525858 159452
rect 176746 159332 176752 159384
rect 176804 159372 176810 159384
rect 258350 159372 258356 159384
rect 176804 159344 258356 159372
rect 176804 159332 176810 159344
rect 258350 159332 258356 159344
rect 258408 159332 258414 159384
rect 285858 159332 285864 159384
rect 285916 159372 285922 159384
rect 529934 159372 529940 159384
rect 285916 159344 529940 159372
rect 285916 159332 285922 159344
rect 529934 159332 529940 159344
rect 529992 159332 529998 159384
rect 255222 158652 255228 158704
rect 255280 158692 255286 158704
rect 269390 158692 269396 158704
rect 255280 158664 269396 158692
rect 255280 158652 255286 158664
rect 269390 158652 269396 158664
rect 269448 158652 269454 158704
rect 272886 158652 272892 158704
rect 272944 158692 272950 158704
rect 300854 158692 300860 158704
rect 272944 158664 300860 158692
rect 272944 158652 272950 158664
rect 300854 158652 300860 158664
rect 300912 158652 300918 158704
rect 301498 158652 301504 158704
rect 301556 158692 301562 158704
rect 345566 158692 345572 158704
rect 301556 158664 345572 158692
rect 301556 158652 301562 158664
rect 345566 158652 345572 158664
rect 345624 158652 345630 158704
rect 249702 158584 249708 158636
rect 249760 158624 249766 158636
rect 265342 158624 265348 158636
rect 249760 158596 265348 158624
rect 249760 158584 249766 158596
rect 265342 158584 265348 158596
rect 265400 158584 265406 158636
rect 272058 158584 272064 158636
rect 272116 158624 272122 158636
rect 346946 158624 346952 158636
rect 272116 158596 346952 158624
rect 272116 158584 272122 158596
rect 346946 158584 346952 158596
rect 347004 158584 347010 158636
rect 251082 158516 251088 158568
rect 251140 158556 251146 158568
rect 266814 158556 266820 158568
rect 251140 158528 266820 158556
rect 251140 158516 251146 158528
rect 266814 158516 266820 158528
rect 266872 158516 266878 158568
rect 271138 158516 271144 158568
rect 271196 158556 271202 158568
rect 348050 158556 348056 158568
rect 271196 158528 348056 158556
rect 271196 158516 271202 158528
rect 348050 158516 348056 158528
rect 348108 158516 348114 158568
rect 249610 158448 249616 158500
rect 249668 158488 249674 158500
rect 267918 158488 267924 158500
rect 249668 158460 267924 158488
rect 249668 158448 249674 158460
rect 267918 158448 267924 158460
rect 267976 158448 267982 158500
rect 272242 158448 272248 158500
rect 272300 158488 272306 158500
rect 349706 158488 349712 158500
rect 272300 158460 349712 158488
rect 272300 158448 272306 158460
rect 349706 158448 349712 158460
rect 349764 158448 349770 158500
rect 246666 158380 246672 158432
rect 246724 158420 246730 158432
rect 266722 158420 266728 158432
rect 246724 158392 266728 158420
rect 246724 158380 246730 158392
rect 266722 158380 266728 158392
rect 266780 158380 266786 158432
rect 270954 158380 270960 158432
rect 271012 158420 271018 158432
rect 349522 158420 349528 158432
rect 271012 158392 349528 158420
rect 271012 158380 271018 158392
rect 349522 158380 349528 158392
rect 349580 158380 349586 158432
rect 246758 158312 246764 158364
rect 246816 158352 246822 158364
rect 246816 158324 263916 158352
rect 246816 158312 246822 158324
rect 242986 158244 242992 158296
rect 243044 158284 243050 158296
rect 263778 158284 263784 158296
rect 243044 158256 263784 158284
rect 243044 158244 243050 158256
rect 263778 158244 263784 158256
rect 263836 158244 263842 158296
rect 263888 158284 263916 158324
rect 264514 158312 264520 158364
rect 264572 158352 264578 158364
rect 265618 158352 265624 158364
rect 264572 158324 265624 158352
rect 264572 158312 264578 158324
rect 265618 158312 265624 158324
rect 265676 158312 265682 158364
rect 271046 158312 271052 158364
rect 271104 158352 271110 158364
rect 349798 158352 349804 158364
rect 271104 158324 349804 158352
rect 271104 158312 271110 158324
rect 349798 158312 349804 158324
rect 349856 158312 349862 158364
rect 266906 158284 266912 158296
rect 263888 158256 266912 158284
rect 266906 158244 266912 158256
rect 266964 158244 266970 158296
rect 269482 158244 269488 158296
rect 269540 158284 269546 158296
rect 349614 158284 349620 158296
rect 269540 158256 349620 158284
rect 269540 158244 269546 158256
rect 349614 158244 349620 158256
rect 349672 158244 349678 158296
rect 219434 158176 219440 158228
rect 219492 158216 219498 158228
rect 262858 158216 262864 158228
rect 219492 158188 262864 158216
rect 219492 158176 219498 158188
rect 262858 158176 262864 158188
rect 262916 158176 262922 158228
rect 272150 158176 272156 158228
rect 272208 158216 272214 158228
rect 353294 158216 353300 158228
rect 272208 158188 353300 158216
rect 272208 158176 272214 158188
rect 353294 158176 353300 158188
rect 353352 158176 353358 158228
rect 208394 158108 208400 158160
rect 208452 158148 208458 158160
rect 261202 158148 261208 158160
rect 208452 158120 261208 158148
rect 208452 158108 208458 158120
rect 261202 158108 261208 158120
rect 261260 158108 261266 158160
rect 271966 158108 271972 158160
rect 272024 158148 272030 158160
rect 357526 158148 357532 158160
rect 272024 158120 357532 158148
rect 272024 158108 272030 158120
rect 357526 158108 357532 158120
rect 357584 158108 357590 158160
rect 204254 158040 204260 158092
rect 204312 158080 204318 158092
rect 261110 158080 261116 158092
rect 204312 158052 261116 158080
rect 204312 158040 204318 158052
rect 261110 158040 261116 158052
rect 261168 158040 261174 158092
rect 284478 158040 284484 158092
rect 284536 158080 284542 158092
rect 284536 158052 291884 158080
rect 284536 158040 284542 158052
rect 187694 157972 187700 158024
rect 187752 158012 187758 158024
rect 259822 158012 259828 158024
rect 187752 157984 259828 158012
rect 187752 157972 187758 157984
rect 259822 157972 259828 157984
rect 259880 157972 259886 158024
rect 259914 157972 259920 158024
rect 259972 158012 259978 158024
rect 260558 158012 260564 158024
rect 259972 157984 260564 158012
rect 259972 157972 259978 157984
rect 260558 157972 260564 157984
rect 260616 157972 260622 158024
rect 281258 157972 281264 158024
rect 281316 158012 281322 158024
rect 287698 158012 287704 158024
rect 281316 157984 287704 158012
rect 281316 157972 281322 157984
rect 287698 157972 287704 157984
rect 287756 157972 287762 158024
rect 291856 158012 291884 158052
rect 293218 158040 293224 158092
rect 293276 158080 293282 158092
rect 411254 158080 411260 158092
rect 293276 158052 411260 158080
rect 293276 158040 293282 158052
rect 411254 158040 411260 158052
rect 411312 158040 411318 158092
rect 505094 158012 505100 158024
rect 291856 157984 505100 158012
rect 505094 157972 505100 157984
rect 505152 157972 505158 158024
rect 253842 157904 253848 157956
rect 253900 157944 253906 157956
rect 266630 157944 266636 157956
rect 253900 157916 266636 157944
rect 253900 157904 253906 157916
rect 266630 157904 266636 157916
rect 266688 157904 266694 157956
rect 301682 157904 301688 157956
rect 301740 157944 301746 157956
rect 331490 157944 331496 157956
rect 301740 157916 331496 157944
rect 301740 157904 301746 157916
rect 331490 157904 331496 157916
rect 331548 157904 331554 157956
rect 337378 157904 337384 157956
rect 337436 157944 337442 157956
rect 339862 157944 339868 157956
rect 337436 157916 339868 157944
rect 337436 157904 337442 157916
rect 339862 157904 339868 157916
rect 339920 157904 339926 157956
rect 300302 157836 300308 157888
rect 300360 157876 300366 157888
rect 319254 157876 319260 157888
rect 300360 157848 319260 157876
rect 300360 157836 300366 157848
rect 319254 157836 319260 157848
rect 319312 157836 319318 157888
rect 256786 157768 256792 157820
rect 256844 157808 256850 157820
rect 261478 157808 261484 157820
rect 256844 157780 261484 157808
rect 256844 157768 256850 157780
rect 261478 157768 261484 157780
rect 261536 157768 261542 157820
rect 301590 157768 301596 157820
rect 301648 157808 301654 157820
rect 314746 157808 314752 157820
rect 301648 157780 314752 157808
rect 301648 157768 301654 157780
rect 314746 157768 314752 157780
rect 314804 157768 314810 157820
rect 259822 157428 259828 157480
rect 259880 157468 259886 157480
rect 265250 157468 265256 157480
rect 259880 157440 265256 157468
rect 259880 157428 259886 157440
rect 265250 157428 265256 157440
rect 265308 157428 265314 157480
rect 3602 157360 3608 157412
rect 3660 157400 3666 157412
rect 293954 157400 293960 157412
rect 3660 157372 293960 157400
rect 3660 157360 3666 157372
rect 293954 157360 293960 157372
rect 294012 157360 294018 157412
rect 264238 157060 264244 157072
rect 258046 157032 264244 157060
rect 250438 156884 250444 156936
rect 250496 156924 250502 156936
rect 258046 156924 258074 157032
rect 264238 157020 264244 157032
rect 264296 157020 264302 157072
rect 264330 156992 264336 157004
rect 250496 156896 258074 156924
rect 258276 156964 264336 156992
rect 250496 156884 250502 156896
rect 240134 156816 240140 156868
rect 240192 156856 240198 156868
rect 258276 156856 258304 156964
rect 264330 156952 264336 156964
rect 264388 156952 264394 157004
rect 300118 156952 300124 157004
rect 300176 156992 300182 157004
rect 345014 156992 345020 157004
rect 300176 156964 345020 156992
rect 300176 156952 300182 156964
rect 345014 156952 345020 156964
rect 345072 156952 345078 157004
rect 300210 156884 300216 156936
rect 300268 156924 300274 156936
rect 345750 156924 345756 156936
rect 300268 156896 345756 156924
rect 300268 156884 300274 156896
rect 345750 156884 345756 156896
rect 345808 156884 345814 156936
rect 262674 156856 262680 156868
rect 240192 156828 258304 156856
rect 258460 156828 262680 156856
rect 240192 156816 240198 156828
rect 231854 156748 231860 156800
rect 231912 156788 231918 156800
rect 258460 156788 258488 156828
rect 262674 156816 262680 156828
rect 262732 156816 262738 156868
rect 273254 156816 273260 156868
rect 273312 156856 273318 156868
rect 360194 156856 360200 156868
rect 273312 156828 360200 156856
rect 273312 156816 273318 156828
rect 360194 156816 360200 156828
rect 360252 156816 360258 156868
rect 261018 156788 261024 156800
rect 231912 156760 258488 156788
rect 258552 156760 261024 156788
rect 231912 156748 231918 156760
rect 213914 156680 213920 156732
rect 213972 156720 213978 156732
rect 258552 156720 258580 156760
rect 261018 156748 261024 156760
rect 261076 156748 261082 156800
rect 281534 156748 281540 156800
rect 281592 156788 281598 156800
rect 473446 156788 473452 156800
rect 281592 156760 473452 156788
rect 281592 156748 281598 156760
rect 473446 156748 473452 156760
rect 473504 156748 473510 156800
rect 213972 156692 258580 156720
rect 213972 156680 213978 156692
rect 259638 156680 259644 156732
rect 259696 156720 259702 156732
rect 265158 156720 265164 156732
rect 259696 156692 265164 156720
rect 259696 156680 259702 156692
rect 265158 156680 265164 156692
rect 265216 156680 265222 156732
rect 283006 156680 283012 156732
rect 283064 156720 283070 156732
rect 495434 156720 495440 156732
rect 283064 156692 495440 156720
rect 283064 156680 283070 156692
rect 495434 156680 495440 156692
rect 495492 156680 495498 156732
rect 205634 156612 205640 156664
rect 205692 156652 205698 156664
rect 205692 156624 258074 156652
rect 205692 156612 205698 156624
rect 258046 156584 258074 156624
rect 259730 156612 259736 156664
rect 259788 156652 259794 156664
rect 260742 156652 260748 156664
rect 259788 156624 260748 156652
rect 259788 156612 259794 156624
rect 260742 156612 260748 156624
rect 260800 156612 260806 156664
rect 285306 156612 285312 156664
rect 285364 156652 285370 156664
rect 502334 156652 502340 156664
rect 285364 156624 502340 156652
rect 285364 156612 285370 156624
rect 502334 156612 502340 156624
rect 502392 156612 502398 156664
rect 261662 156584 261668 156596
rect 258046 156556 261668 156584
rect 261662 156544 261668 156556
rect 261720 156544 261726 156596
rect 259914 156000 259920 156052
rect 259972 156040 259978 156052
rect 260374 156040 260380 156052
rect 259972 156012 260380 156040
rect 259972 156000 259978 156012
rect 260374 156000 260380 156012
rect 260432 156000 260438 156052
rect 259270 155864 259276 155916
rect 259328 155904 259334 155916
rect 265526 155904 265532 155916
rect 259328 155876 265532 155904
rect 259328 155864 259334 155876
rect 265526 155864 265532 155876
rect 265584 155864 265590 155916
rect 259086 155796 259092 155848
rect 259144 155836 259150 155848
rect 266538 155836 266544 155848
rect 259144 155808 266544 155836
rect 259144 155796 259150 155808
rect 266538 155796 266544 155808
rect 266596 155796 266602 155848
rect 270862 155796 270868 155848
rect 270920 155836 270926 155848
rect 270920 155808 277394 155836
rect 270920 155796 270926 155808
rect 259178 155728 259184 155780
rect 259236 155768 259242 155780
rect 267550 155768 267556 155780
rect 259236 155740 267556 155768
rect 259236 155728 259242 155740
rect 267550 155728 267556 155740
rect 267608 155728 267614 155780
rect 270770 155728 270776 155780
rect 270828 155768 270834 155780
rect 270828 155740 272012 155768
rect 270828 155728 270834 155740
rect 260282 155660 260288 155712
rect 260340 155700 260346 155712
rect 261570 155700 261576 155712
rect 260340 155672 261576 155700
rect 260340 155660 260346 155672
rect 261570 155660 261576 155672
rect 261628 155660 261634 155712
rect 270678 155660 270684 155712
rect 270736 155700 270742 155712
rect 271874 155700 271880 155712
rect 270736 155672 271880 155700
rect 270736 155660 270742 155672
rect 271874 155660 271880 155672
rect 271932 155660 271938 155712
rect 257706 155592 257712 155644
rect 257764 155632 257770 155644
rect 267826 155632 267832 155644
rect 257764 155604 267832 155632
rect 257764 155592 257770 155604
rect 267826 155592 267832 155604
rect 267884 155592 267890 155644
rect 269114 155592 269120 155644
rect 269172 155632 269178 155644
rect 269172 155604 271828 155632
rect 269172 155592 269178 155604
rect 257522 155524 257528 155576
rect 257580 155564 257586 155576
rect 268654 155564 268660 155576
rect 257580 155536 268660 155564
rect 257580 155524 257586 155536
rect 268654 155524 268660 155536
rect 268712 155524 268718 155576
rect 253750 155456 253756 155508
rect 253808 155496 253814 155508
rect 265802 155496 265808 155508
rect 253808 155468 265808 155496
rect 253808 155456 253814 155468
rect 265802 155456 265808 155468
rect 265860 155456 265866 155508
rect 197354 155388 197360 155440
rect 197412 155428 197418 155440
rect 260006 155428 260012 155440
rect 197412 155400 260012 155428
rect 197412 155388 197418 155400
rect 260006 155388 260012 155400
rect 260064 155388 260070 155440
rect 260466 155388 260472 155440
rect 260524 155388 260530 155440
rect 270586 155388 270592 155440
rect 270644 155428 270650 155440
rect 271690 155428 271696 155440
rect 270644 155400 270816 155428
rect 270644 155388 270650 155400
rect 194594 155320 194600 155372
rect 194652 155360 194658 155372
rect 259454 155360 259460 155372
rect 194652 155332 259460 155360
rect 194652 155320 194658 155332
rect 259454 155320 259460 155332
rect 259512 155320 259518 155372
rect 193306 155252 193312 155304
rect 193364 155292 193370 155304
rect 260484 155292 260512 155388
rect 193364 155264 260512 155292
rect 193364 155252 193370 155264
rect 190454 155184 190460 155236
rect 190512 155224 190518 155236
rect 259914 155224 259920 155236
rect 190512 155196 259920 155224
rect 190512 155184 190518 155196
rect 259914 155184 259920 155196
rect 259972 155184 259978 155236
rect 270788 155224 270816 155400
rect 271524 155400 271696 155428
rect 271524 155292 271552 155400
rect 271690 155388 271696 155400
rect 271748 155388 271754 155440
rect 271800 155360 271828 155604
rect 271984 155496 272012 155740
rect 277366 155564 277394 155808
rect 344186 155564 344192 155576
rect 277366 155536 344192 155564
rect 344186 155524 344192 155536
rect 344244 155524 344250 155576
rect 344370 155496 344376 155508
rect 271984 155468 344376 155496
rect 344370 155456 344376 155468
rect 344428 155456 344434 155508
rect 271874 155388 271880 155440
rect 271932 155428 271938 155440
rect 344462 155428 344468 155440
rect 271932 155400 344468 155428
rect 271932 155388 271938 155400
rect 344462 155388 344468 155400
rect 344520 155388 344526 155440
rect 344554 155360 344560 155372
rect 271800 155332 344560 155360
rect 344554 155320 344560 155332
rect 344612 155320 344618 155372
rect 347130 155292 347136 155304
rect 271524 155264 347136 155292
rect 347130 155252 347136 155264
rect 347188 155252 347194 155304
rect 347222 155224 347228 155236
rect 270788 155196 347228 155224
rect 347222 155184 347228 155196
rect 347280 155184 347286 155236
rect 30374 153824 30380 153876
rect 30432 153864 30438 153876
rect 247494 153864 247500 153876
rect 30432 153836 247500 153864
rect 30432 153824 30438 153836
rect 247494 153824 247500 153836
rect 247552 153824 247558 153876
rect 233970 153144 233976 153196
rect 234028 153184 234034 153196
rect 256694 153184 256700 153196
rect 234028 153156 256700 153184
rect 234028 153144 234034 153156
rect 256694 153144 256700 153156
rect 256752 153144 256758 153196
rect 3326 150356 3332 150408
rect 3384 150396 3390 150408
rect 94498 150396 94504 150408
rect 3384 150368 94504 150396
rect 3384 150356 3390 150368
rect 94498 150356 94504 150368
rect 94556 150356 94562 150408
rect 234154 144848 234160 144900
rect 234212 144888 234218 144900
rect 256694 144888 256700 144900
rect 234212 144860 256700 144888
rect 234212 144848 234218 144860
rect 256694 144848 256700 144860
rect 256752 144848 256758 144900
rect 257246 142060 257252 142112
rect 257304 142100 257310 142112
rect 257798 142100 257804 142112
rect 257304 142072 257804 142100
rect 257304 142060 257310 142072
rect 257798 142060 257804 142072
rect 257856 142060 257862 142112
rect 577682 139340 577688 139392
rect 577740 139380 577746 139392
rect 579614 139380 579620 139392
rect 577740 139352 579620 139380
rect 577740 139340 577746 139352
rect 579614 139340 579620 139352
rect 579672 139340 579678 139392
rect 3050 137912 3056 137964
rect 3108 137952 3114 137964
rect 235258 137952 235264 137964
rect 3108 137924 235264 137952
rect 3108 137912 3114 137924
rect 235258 137912 235264 137924
rect 235316 137912 235322 137964
rect 234246 135192 234252 135244
rect 234304 135232 234310 135244
rect 256786 135232 256792 135244
rect 234304 135204 256792 135232
rect 234304 135192 234310 135204
rect 256786 135192 256792 135204
rect 256844 135192 256850 135244
rect 232498 131044 232504 131096
rect 232556 131084 232562 131096
rect 256786 131084 256792 131096
rect 232556 131056 256792 131084
rect 232556 131044 232562 131056
rect 256786 131044 256792 131056
rect 256844 131044 256850 131096
rect 344278 130364 344284 130416
rect 344336 130404 344342 130416
rect 345014 130404 345020 130416
rect 344336 130376 345020 130404
rect 344336 130364 344342 130376
rect 345014 130364 345020 130376
rect 345072 130364 345078 130416
rect 234798 126896 234804 126948
rect 234856 126936 234862 126948
rect 235626 126936 235632 126948
rect 234856 126908 235632 126936
rect 234856 126896 234862 126908
rect 235626 126896 235632 126908
rect 235684 126936 235690 126948
rect 256786 126936 256792 126948
rect 235684 126908 256792 126936
rect 235684 126896 235690 126908
rect 256786 126896 256792 126908
rect 256844 126896 256850 126948
rect 347038 126896 347044 126948
rect 347096 126936 347102 126948
rect 579706 126936 579712 126948
rect 347096 126908 579712 126936
rect 347096 126896 347102 126908
rect 579706 126896 579712 126908
rect 579764 126896 579770 126948
rect 90450 126216 90456 126268
rect 90508 126256 90514 126268
rect 234798 126256 234804 126268
rect 90508 126228 234804 126256
rect 90508 126216 90514 126228
rect 234798 126216 234804 126228
rect 234856 126216 234862 126268
rect 235718 122748 235724 122800
rect 235776 122788 235782 122800
rect 256786 122788 256792 122800
rect 235776 122760 256792 122788
rect 235776 122748 235782 122760
rect 256786 122748 256792 122760
rect 256844 122748 256850 122800
rect 234338 113092 234344 113144
rect 234396 113132 234402 113144
rect 256786 113132 256792 113144
rect 234396 113104 256792 113132
rect 234396 113092 234402 113104
rect 256786 113092 256792 113104
rect 256844 113092 256850 113144
rect 234522 104796 234528 104848
rect 234580 104836 234586 104848
rect 256786 104836 256792 104848
rect 234580 104808 256792 104836
rect 234580 104796 234586 104808
rect 256786 104796 256792 104808
rect 256844 104796 256850 104848
rect 577590 100648 577596 100700
rect 577648 100688 577654 100700
rect 579614 100688 579620 100700
rect 577648 100660 579620 100688
rect 577648 100648 577654 100660
rect 579614 100648 579620 100660
rect 579672 100648 579678 100700
rect 259730 100444 259736 100496
rect 259788 100484 259794 100496
rect 263686 100484 263692 100496
rect 259788 100456 263692 100484
rect 259788 100444 259794 100456
rect 263686 100444 263692 100456
rect 263744 100444 263750 100496
rect 256510 100036 256516 100088
rect 256568 100076 256574 100088
rect 260834 100076 260840 100088
rect 256568 100048 260840 100076
rect 256568 100036 256574 100048
rect 260834 100036 260840 100048
rect 260892 100036 260898 100088
rect 246942 99968 246948 100020
rect 247000 100008 247006 100020
rect 262214 100008 262220 100020
rect 247000 99980 262220 100008
rect 247000 99968 247006 99980
rect 262214 99968 262220 99980
rect 262272 99968 262278 100020
rect 257982 97928 257988 97980
rect 258040 97968 258046 97980
rect 267734 97968 267740 97980
rect 258040 97940 267740 97968
rect 258040 97928 258046 97940
rect 267734 97928 267740 97940
rect 267792 97928 267798 97980
rect 334710 97928 334716 97980
rect 334768 97968 334774 97980
rect 349890 97968 349896 97980
rect 334768 97940 349896 97968
rect 334768 97928 334774 97940
rect 349890 97928 349896 97940
rect 349948 97928 349954 97980
rect 245102 97860 245108 97912
rect 245160 97900 245166 97912
rect 297358 97900 297364 97912
rect 245160 97872 297364 97900
rect 245160 97860 245166 97872
rect 297358 97860 297364 97872
rect 297416 97860 297422 97912
rect 317966 97860 317972 97912
rect 318024 97900 318030 97912
rect 349246 97900 349252 97912
rect 318024 97872 349252 97900
rect 318024 97860 318030 97872
rect 349246 97860 349252 97872
rect 349304 97860 349310 97912
rect 258994 97792 259000 97844
rect 259052 97832 259058 97844
rect 301222 97832 301228 97844
rect 259052 97804 301228 97832
rect 259052 97792 259058 97804
rect 301222 97792 301228 97804
rect 301280 97792 301286 97844
rect 339218 97792 339224 97844
rect 339276 97832 339282 97844
rect 347866 97832 347872 97844
rect 339276 97804 347872 97832
rect 339276 97792 339282 97804
rect 347866 97792 347872 97804
rect 347924 97792 347930 97844
rect 257890 97724 257896 97776
rect 257948 97764 257954 97776
rect 276106 97764 276112 97776
rect 257948 97736 276112 97764
rect 257948 97724 257954 97736
rect 276106 97724 276112 97736
rect 276164 97724 276170 97776
rect 322474 97724 322480 97776
rect 322532 97764 322538 97776
rect 347774 97764 347780 97776
rect 322532 97736 347780 97764
rect 322532 97724 322538 97736
rect 347774 97724 347780 97736
rect 347832 97724 347838 97776
rect 259546 97656 259552 97708
rect 259604 97696 259610 97708
rect 284478 97696 284484 97708
rect 259604 97668 284484 97696
rect 259604 97656 259610 97668
rect 284478 97656 284484 97668
rect 284536 97656 284542 97708
rect 326338 97656 326344 97708
rect 326396 97696 326402 97708
rect 348326 97696 348332 97708
rect 326396 97668 348332 97696
rect 326396 97656 326402 97668
rect 348326 97656 348332 97668
rect 348384 97656 348390 97708
rect 257338 97588 257344 97640
rect 257396 97628 257402 97640
rect 280614 97628 280620 97640
rect 257396 97600 280620 97628
rect 257396 97588 257402 97600
rect 280614 97588 280620 97600
rect 280672 97588 280678 97640
rect 309594 97588 309600 97640
rect 309652 97628 309658 97640
rect 344646 97628 344652 97640
rect 309652 97600 344652 97628
rect 309652 97588 309658 97600
rect 344646 97588 344652 97600
rect 344704 97588 344710 97640
rect 234430 97520 234436 97572
rect 234488 97560 234494 97572
rect 292850 97560 292856 97572
rect 234488 97532 292856 97560
rect 234488 97520 234494 97532
rect 292850 97520 292856 97532
rect 292908 97520 292914 97572
rect 314102 97520 314108 97572
rect 314160 97560 314166 97572
rect 344002 97560 344008 97572
rect 314160 97532 344008 97560
rect 314160 97520 314166 97532
rect 344002 97520 344008 97532
rect 344060 97520 344066 97572
rect 235810 97452 235816 97504
rect 235868 97492 235874 97504
rect 263870 97492 263876 97504
rect 235868 97464 263876 97492
rect 235868 97452 235874 97464
rect 263870 97452 263876 97464
rect 263928 97452 263934 97504
rect 99374 89020 99380 89072
rect 99432 89060 99438 89072
rect 243814 89060 243820 89072
rect 99432 89032 243820 89060
rect 99432 89020 99438 89032
rect 243814 89020 243820 89032
rect 243872 89020 243878 89072
rect 92474 88952 92480 89004
rect 92532 88992 92538 89004
rect 243906 88992 243912 89004
rect 92532 88964 243912 88992
rect 92532 88952 92538 88964
rect 243906 88952 243912 88964
rect 243964 88952 243970 89004
rect 3326 85484 3332 85536
rect 3384 85524 3390 85536
rect 90358 85524 90364 85536
rect 3384 85496 90364 85524
rect 3384 85484 3390 85496
rect 90358 85484 90364 85496
rect 90416 85484 90422 85536
rect 86954 82084 86960 82136
rect 87012 82124 87018 82136
rect 251542 82124 251548 82136
rect 87012 82096 251548 82124
rect 87012 82084 87018 82096
rect 251542 82084 251548 82096
rect 251600 82084 251606 82136
rect 3326 71680 3332 71732
rect 3384 71720 3390 71732
rect 235902 71720 235908 71732
rect 3384 71692 235908 71720
rect 3384 71680 3390 71692
rect 235902 71680 235908 71692
rect 235960 71720 235966 71732
rect 304994 71720 305000 71732
rect 235960 71692 305000 71720
rect 235960 71680 235966 71692
rect 304994 71680 305000 71692
rect 305052 71680 305058 71732
rect 3326 59304 3332 59356
rect 3384 59344 3390 59356
rect 231118 59344 231124 59356
rect 3384 59316 231124 59344
rect 3384 59304 3390 59316
rect 231118 59304 231124 59316
rect 231176 59304 231182 59356
rect 3510 33056 3516 33108
rect 3568 33096 3574 33108
rect 90450 33096 90456 33108
rect 3568 33068 90456 33096
rect 3568 33056 3574 33068
rect 90450 33056 90456 33068
rect 90508 33056 90514 33108
rect 142154 21360 142160 21412
rect 142212 21400 142218 21412
rect 255590 21400 255596 21412
rect 142212 21372 255596 21400
rect 142212 21360 142218 21372
rect 255590 21360 255596 21372
rect 255648 21360 255654 21412
rect 3510 20612 3516 20664
rect 3568 20652 3574 20664
rect 174538 20652 174544 20664
rect 3568 20624 174544 20652
rect 3568 20612 3574 20624
rect 174538 20612 174544 20624
rect 174596 20612 174602 20664
rect 577498 20612 577504 20664
rect 577556 20652 577562 20664
rect 579706 20652 579712 20664
rect 577556 20624 579712 20652
rect 577556 20612 577562 20624
rect 579706 20612 579712 20624
rect 579764 20612 579770 20664
rect 120626 14560 120632 14612
rect 120684 14600 120690 14612
rect 254302 14600 254308 14612
rect 120684 14572 254308 14600
rect 120684 14560 120690 14572
rect 254302 14560 254308 14572
rect 254360 14560 254366 14612
rect 110506 14492 110512 14544
rect 110564 14532 110570 14544
rect 253014 14532 253020 14544
rect 110564 14504 253020 14532
rect 110564 14492 110570 14504
rect 253014 14492 253020 14504
rect 253072 14492 253078 14544
rect 102226 14424 102232 14476
rect 102284 14464 102290 14476
rect 252922 14464 252928 14476
rect 102284 14436 252928 14464
rect 102284 14424 102290 14436
rect 252922 14424 252928 14436
rect 252980 14424 252986 14476
rect 124674 13200 124680 13252
rect 124732 13240 124738 13252
rect 245010 13240 245016 13252
rect 124732 13212 245016 13240
rect 124732 13200 124738 13212
rect 245010 13200 245016 13212
rect 245068 13200 245074 13252
rect 122282 13132 122288 13184
rect 122340 13172 122346 13184
rect 254210 13172 254216 13184
rect 122340 13144 254216 13172
rect 122340 13132 122346 13144
rect 254210 13132 254216 13144
rect 254268 13132 254274 13184
rect 13538 13064 13544 13116
rect 13596 13104 13602 13116
rect 246022 13104 246028 13116
rect 13596 13076 246028 13104
rect 13596 13064 13602 13076
rect 246022 13064 246028 13076
rect 246080 13064 246086 13116
rect 127618 12248 127624 12300
rect 127676 12288 127682 12300
rect 250346 12288 250352 12300
rect 127676 12260 250352 12288
rect 127676 12248 127682 12260
rect 250346 12248 250352 12260
rect 250404 12248 250410 12300
rect 117314 12180 117320 12232
rect 117372 12220 117378 12232
rect 254118 12220 254124 12232
rect 117372 12192 254124 12220
rect 117372 12180 117378 12192
rect 254118 12180 254124 12192
rect 254176 12180 254182 12232
rect 108114 12112 108120 12164
rect 108172 12152 108178 12164
rect 252646 12152 252652 12164
rect 108172 12124 252652 12152
rect 108172 12112 108178 12124
rect 252646 12112 252652 12124
rect 252704 12112 252710 12164
rect 104066 12044 104072 12096
rect 104124 12084 104130 12096
rect 252830 12084 252836 12096
rect 104124 12056 252836 12084
rect 104124 12044 104130 12056
rect 252830 12044 252836 12056
rect 252888 12044 252894 12096
rect 100754 11976 100760 12028
rect 100812 12016 100818 12028
rect 252738 12016 252744 12028
rect 100812 11988 252744 12016
rect 100812 11976 100818 11988
rect 252738 11976 252744 11988
rect 252796 11976 252802 12028
rect 89898 11908 89904 11960
rect 89956 11948 89962 11960
rect 251450 11948 251456 11960
rect 89956 11920 251456 11948
rect 89956 11908 89962 11920
rect 251450 11908 251456 11920
rect 251508 11908 251514 11960
rect 5258 11840 5264 11892
rect 5316 11880 5322 11892
rect 178862 11880 178868 11892
rect 5316 11852 178868 11880
rect 5316 11840 5322 11852
rect 178862 11840 178868 11852
rect 178920 11840 178926 11892
rect 347958 11840 347964 11892
rect 348016 11840 348022 11892
rect 73338 11772 73344 11824
rect 73396 11812 73402 11824
rect 250254 11812 250260 11824
rect 73396 11784 250260 11812
rect 73396 11772 73402 11784
rect 250254 11772 250260 11784
rect 250312 11772 250318 11824
rect 33594 11704 33600 11756
rect 33652 11744 33658 11756
rect 247402 11744 247408 11756
rect 33652 11716 247408 11744
rect 33652 11704 33658 11716
rect 247402 11704 247408 11716
rect 247460 11704 247466 11756
rect 160094 11636 160100 11688
rect 160152 11676 160158 11688
rect 161290 11676 161296 11688
rect 160152 11648 161296 11676
rect 160152 11636 160158 11648
rect 161290 11636 161296 11648
rect 161348 11636 161354 11688
rect 184934 11636 184940 11688
rect 184992 11676 184998 11688
rect 186130 11676 186136 11688
rect 184992 11648 186136 11676
rect 184992 11636 184998 11648
rect 186130 11636 186136 11648
rect 186188 11636 186194 11688
rect 201494 11636 201500 11688
rect 201552 11676 201558 11688
rect 202690 11676 202696 11688
rect 201552 11648 202696 11676
rect 201552 11636 201558 11648
rect 202690 11636 202696 11648
rect 202748 11636 202754 11688
rect 234614 11636 234620 11688
rect 234672 11676 234678 11688
rect 235810 11676 235816 11688
rect 234672 11648 235816 11676
rect 234672 11636 234678 11648
rect 235810 11636 235816 11648
rect 235868 11636 235874 11688
rect 347976 11676 348004 11840
rect 348050 11676 348056 11688
rect 347976 11648 348056 11676
rect 348050 11636 348056 11648
rect 348108 11636 348114 11688
rect 181438 10684 181444 10736
rect 181496 10724 181502 10736
rect 251358 10724 251364 10736
rect 181496 10696 251364 10724
rect 181496 10684 181502 10696
rect 251358 10684 251364 10696
rect 251416 10684 251422 10736
rect 114002 10616 114008 10668
rect 114060 10656 114066 10668
rect 242526 10656 242532 10668
rect 114060 10628 242532 10656
rect 114060 10616 114066 10628
rect 242526 10616 242532 10628
rect 242584 10616 242590 10668
rect 42794 10548 42800 10600
rect 42852 10588 42858 10600
rect 200758 10588 200764 10600
rect 42852 10560 200764 10588
rect 42852 10548 42858 10560
rect 200758 10548 200764 10560
rect 200816 10548 200822 10600
rect 20162 10480 20168 10532
rect 20220 10520 20226 10532
rect 182818 10520 182824 10532
rect 20220 10492 182824 10520
rect 20220 10480 20226 10492
rect 182818 10480 182824 10492
rect 182876 10480 182882 10532
rect 221458 10480 221464 10532
rect 221516 10520 221522 10532
rect 247218 10520 247224 10532
rect 221516 10492 247224 10520
rect 221516 10480 221522 10492
rect 247218 10480 247224 10492
rect 247276 10480 247282 10532
rect 69106 10412 69112 10464
rect 69164 10452 69170 10464
rect 250162 10452 250168 10464
rect 69164 10424 250168 10452
rect 69164 10412 69170 10424
rect 250162 10412 250168 10424
rect 250220 10412 250226 10464
rect 36722 10344 36728 10396
rect 36780 10384 36786 10396
rect 247310 10384 247316 10396
rect 36780 10356 247316 10384
rect 36780 10344 36786 10356
rect 247310 10344 247316 10356
rect 247368 10344 247374 10396
rect 11882 10276 11888 10328
rect 11940 10316 11946 10328
rect 245930 10316 245936 10328
rect 11940 10288 245936 10316
rect 11940 10276 11946 10288
rect 245930 10276 245936 10288
rect 245988 10276 245994 10328
rect 239674 9596 239680 9648
rect 239732 9636 239738 9648
rect 291378 9636 291384 9648
rect 239732 9608 291384 9636
rect 239732 9596 239738 9608
rect 291378 9596 291384 9608
rect 291436 9596 291442 9648
rect 196066 9528 196072 9580
rect 196124 9568 196130 9580
rect 250070 9568 250076 9580
rect 196124 9540 250076 9568
rect 196124 9528 196130 9540
rect 250070 9528 250076 9540
rect 250128 9528 250134 9580
rect 239766 9460 239772 9512
rect 239824 9500 239830 9512
rect 294874 9500 294880 9512
rect 239824 9472 294880 9500
rect 239824 9460 239830 9472
rect 294874 9460 294880 9472
rect 294932 9460 294938 9512
rect 239950 9392 239956 9444
rect 240008 9432 240014 9444
rect 298462 9432 298468 9444
rect 240008 9404 298468 9432
rect 240008 9392 240014 9404
rect 298462 9392 298468 9404
rect 298520 9392 298526 9444
rect 241330 9324 241336 9376
rect 241388 9364 241394 9376
rect 301958 9364 301964 9376
rect 241388 9336 301964 9364
rect 241388 9324 241394 9336
rect 301958 9324 301964 9336
rect 302016 9324 302022 9376
rect 239582 9256 239588 9308
rect 239640 9296 239646 9308
rect 305546 9296 305552 9308
rect 239640 9268 305552 9296
rect 239640 9256 239646 9268
rect 305546 9256 305552 9268
rect 305604 9256 305610 9308
rect 241238 9188 241244 9240
rect 241296 9228 241302 9240
rect 309042 9228 309048 9240
rect 241296 9200 309048 9228
rect 241296 9188 241302 9200
rect 309042 9188 309048 9200
rect 309100 9188 309106 9240
rect 239858 9120 239864 9172
rect 239916 9160 239922 9172
rect 312630 9160 312636 9172
rect 239916 9132 312636 9160
rect 239916 9120 239922 9132
rect 312630 9120 312636 9132
rect 312688 9120 312694 9172
rect 138842 9052 138848 9104
rect 138900 9092 138906 9104
rect 251818 9092 251824 9104
rect 138900 9064 251824 9092
rect 138900 9052 138906 9064
rect 251818 9052 251824 9064
rect 251876 9052 251882 9104
rect 106918 8984 106924 9036
rect 106976 9024 106982 9036
rect 242434 9024 242440 9036
rect 106976 8996 242440 9024
rect 106976 8984 106982 8996
rect 242434 8984 242440 8996
rect 242492 8984 242498 9036
rect 243998 8984 244004 9036
rect 244056 9024 244062 9036
rect 287790 9024 287796 9036
rect 244056 8996 287796 9024
rect 244056 8984 244062 8996
rect 287790 8984 287796 8996
rect 287848 8984 287854 9036
rect 35986 8916 35992 8968
rect 36044 8956 36050 8968
rect 196618 8956 196624 8968
rect 36044 8928 196624 8956
rect 36044 8916 36050 8928
rect 196618 8916 196624 8928
rect 196676 8916 196682 8968
rect 241146 8916 241152 8968
rect 241204 8956 241210 8968
rect 316218 8956 316224 8968
rect 241204 8928 316224 8956
rect 241204 8916 241210 8928
rect 316218 8916 316224 8928
rect 316276 8916 316282 8968
rect 240042 8848 240048 8900
rect 240100 8888 240106 8900
rect 284294 8888 284300 8900
rect 240100 8860 284300 8888
rect 240100 8848 240106 8860
rect 284294 8848 284300 8860
rect 284352 8848 284358 8900
rect 242066 8780 242072 8832
rect 242124 8820 242130 8832
rect 280706 8820 280712 8832
rect 242124 8792 280712 8820
rect 242124 8780 242130 8792
rect 280706 8780 280712 8792
rect 280764 8780 280770 8832
rect 242618 8712 242624 8764
rect 242676 8752 242682 8764
rect 277118 8752 277124 8764
rect 242676 8724 277124 8752
rect 242676 8712 242682 8724
rect 277118 8712 277124 8724
rect 277176 8712 277182 8764
rect 170766 8032 170772 8084
rect 170824 8072 170830 8084
rect 258718 8072 258724 8084
rect 170824 8044 258724 8072
rect 170824 8032 170830 8044
rect 258718 8032 258724 8044
rect 258776 8032 258782 8084
rect 143534 7964 143540 8016
rect 143592 8004 143598 8016
rect 255498 8004 255504 8016
rect 143592 7976 255504 8004
rect 143592 7964 143598 7976
rect 255498 7964 255504 7976
rect 255556 7964 255562 8016
rect 103330 7896 103336 7948
rect 103388 7936 103394 7948
rect 253658 7936 253664 7948
rect 103388 7908 253664 7936
rect 103388 7896 103394 7908
rect 253658 7896 253664 7908
rect 253716 7896 253722 7948
rect 85666 7828 85672 7880
rect 85724 7868 85730 7880
rect 243722 7868 243728 7880
rect 85724 7840 243728 7868
rect 85724 7828 85730 7840
rect 243722 7828 243728 7840
rect 243780 7828 243786 7880
rect 28902 7760 28908 7812
rect 28960 7800 28966 7812
rect 188338 7800 188344 7812
rect 28960 7772 188344 7800
rect 28960 7760 28966 7772
rect 188338 7760 188344 7772
rect 188396 7760 188402 7812
rect 199102 7760 199108 7812
rect 199160 7800 199166 7812
rect 254578 7800 254584 7812
rect 199160 7772 254584 7800
rect 199160 7760 199166 7772
rect 254578 7760 254584 7772
rect 254636 7760 254642 7812
rect 11146 7692 11152 7744
rect 11204 7732 11210 7744
rect 178678 7732 178684 7744
rect 11204 7704 178684 7732
rect 11204 7692 11210 7704
rect 178678 7692 178684 7704
rect 178736 7692 178742 7744
rect 180242 7692 180248 7744
rect 180300 7732 180306 7744
rect 258258 7732 258264 7744
rect 180300 7704 258264 7732
rect 180300 7692 180306 7704
rect 258258 7692 258264 7704
rect 258316 7692 258322 7744
rect 83274 7624 83280 7676
rect 83332 7664 83338 7676
rect 252094 7664 252100 7676
rect 83332 7636 252100 7664
rect 83332 7624 83338 7636
rect 252094 7624 252100 7636
rect 252152 7624 252158 7676
rect 51350 7556 51356 7608
rect 51408 7596 51414 7608
rect 249518 7596 249524 7608
rect 51408 7568 249524 7596
rect 51408 7556 51414 7568
rect 249518 7556 249524 7568
rect 249576 7556 249582 7608
rect 246758 6808 246764 6860
rect 246816 6848 246822 6860
rect 279510 6848 279516 6860
rect 246816 6820 279516 6848
rect 246816 6808 246822 6820
rect 279510 6808 279516 6820
rect 279568 6808 279574 6860
rect 344922 6808 344928 6860
rect 344980 6848 344986 6860
rect 580166 6848 580172 6860
rect 344980 6820 580172 6848
rect 344980 6808 344986 6820
rect 580166 6808 580172 6820
rect 580224 6808 580230 6860
rect 246666 6740 246672 6792
rect 246724 6780 246730 6792
rect 283098 6780 283104 6792
rect 246724 6752 283104 6780
rect 246724 6740 246730 6752
rect 283098 6740 283104 6752
rect 283156 6740 283162 6792
rect 248322 6672 248328 6724
rect 248380 6712 248386 6724
rect 286594 6712 286600 6724
rect 248380 6684 286600 6712
rect 248380 6672 248386 6684
rect 286594 6672 286600 6684
rect 286652 6672 286658 6724
rect 244090 6604 244096 6656
rect 244148 6644 244154 6656
rect 293678 6644 293684 6656
rect 244148 6616 293684 6644
rect 244148 6604 244154 6616
rect 293678 6604 293684 6616
rect 293736 6604 293742 6656
rect 246850 6536 246856 6588
rect 246908 6576 246914 6588
rect 300762 6576 300768 6588
rect 246908 6548 300768 6576
rect 246908 6536 246914 6548
rect 300762 6536 300768 6548
rect 300820 6536 300826 6588
rect 248230 6468 248236 6520
rect 248288 6508 248294 6520
rect 304350 6508 304356 6520
rect 248288 6480 304356 6508
rect 248288 6468 248294 6480
rect 304350 6468 304356 6480
rect 304408 6468 304414 6520
rect 245470 6400 245476 6452
rect 245528 6440 245534 6452
rect 307938 6440 307944 6452
rect 245528 6412 307944 6440
rect 245528 6400 245534 6412
rect 307938 6400 307944 6412
rect 307996 6400 308002 6452
rect 173158 6332 173164 6384
rect 173216 6372 173222 6384
rect 258534 6372 258540 6384
rect 173216 6344 258540 6372
rect 173216 6332 173222 6344
rect 258534 6332 258540 6344
rect 258592 6332 258598 6384
rect 78582 6264 78588 6316
rect 78640 6304 78646 6316
rect 249150 6304 249156 6316
rect 78640 6276 249156 6304
rect 78640 6264 78646 6276
rect 249150 6264 249156 6276
rect 249208 6264 249214 6316
rect 249610 6264 249616 6316
rect 249668 6304 249674 6316
rect 290182 6304 290188 6316
rect 249668 6276 290188 6304
rect 249668 6264 249674 6276
rect 290182 6264 290188 6276
rect 290240 6264 290246 6316
rect 72602 6196 72608 6248
rect 72660 6236 72666 6248
rect 249978 6236 249984 6248
rect 72660 6208 249984 6236
rect 72660 6196 72666 6208
rect 249978 6196 249984 6208
rect 250036 6196 250042 6248
rect 250990 6196 250996 6248
rect 251048 6236 251054 6248
rect 297266 6236 297272 6248
rect 251048 6208 297272 6236
rect 251048 6196 251054 6208
rect 297266 6196 297272 6208
rect 297324 6196 297330 6248
rect 337470 6196 337476 6248
rect 337528 6236 337534 6248
rect 348234 6236 348240 6248
rect 337528 6208 348240 6236
rect 337528 6196 337534 6208
rect 348234 6196 348240 6208
rect 348292 6196 348298 6248
rect 19426 6128 19432 6180
rect 19484 6168 19490 6180
rect 242342 6168 242348 6180
rect 19484 6140 242348 6168
rect 19484 6128 19490 6140
rect 242342 6128 242348 6140
rect 242400 6128 242406 6180
rect 245562 6128 245568 6180
rect 245620 6168 245626 6180
rect 311434 6168 311440 6180
rect 245620 6140 311440 6168
rect 245620 6128 245626 6140
rect 311434 6128 311440 6140
rect 311492 6128 311498 6180
rect 333882 6128 333888 6180
rect 333940 6168 333946 6180
rect 349798 6168 349804 6180
rect 333940 6140 349804 6168
rect 333940 6128 333946 6140
rect 349798 6128 349804 6140
rect 349856 6128 349862 6180
rect 242710 6060 242716 6112
rect 242768 6100 242774 6112
rect 273622 6100 273628 6112
rect 242768 6072 273628 6100
rect 242768 6060 242774 6072
rect 273622 6060 273628 6072
rect 273680 6060 273686 6112
rect 241422 5992 241428 6044
rect 241480 6032 241486 6044
rect 270034 6032 270040 6044
rect 241480 6004 270040 6032
rect 241480 5992 241486 6004
rect 270034 5992 270040 6004
rect 270092 5992 270098 6044
rect 242802 5924 242808 5976
rect 242860 5964 242866 5976
rect 266538 5964 266544 5976
rect 242860 5936 266544 5964
rect 242860 5924 242866 5936
rect 266538 5924 266544 5936
rect 266596 5924 266602 5976
rect 197354 5108 197360 5160
rect 197412 5148 197418 5160
rect 255774 5148 255780 5160
rect 197412 5120 255780 5148
rect 197412 5108 197418 5120
rect 255774 5108 255780 5120
rect 255832 5108 255838 5160
rect 175918 5040 175924 5092
rect 175976 5080 175982 5092
rect 244274 5080 244280 5092
rect 175976 5052 244280 5080
rect 175976 5040 175982 5052
rect 244274 5040 244280 5052
rect 244332 5040 244338 5092
rect 64322 4972 64328 5024
rect 64380 5012 64386 5024
rect 250806 5012 250812 5024
rect 64380 4984 250812 5012
rect 64380 4972 64386 4984
rect 250806 4972 250812 4984
rect 250864 4972 250870 5024
rect 57238 4904 57244 4956
rect 57296 4944 57302 4956
rect 248966 4944 248972 4956
rect 57296 4916 248972 4944
rect 57296 4904 57302 4916
rect 248966 4904 248972 4916
rect 249024 4904 249030 4956
rect 14734 4836 14740 4888
rect 14792 4876 14798 4888
rect 246206 4876 246212 4888
rect 14792 4848 246212 4876
rect 14792 4836 14798 4848
rect 246206 4836 246212 4848
rect 246264 4836 246270 4888
rect 1670 4768 1676 4820
rect 1728 4808 1734 4820
rect 244366 4808 244372 4820
rect 1728 4780 244372 4808
rect 1728 4768 1734 4780
rect 244366 4768 244372 4780
rect 244424 4768 244430 4820
rect 253842 4088 253848 4140
rect 253900 4128 253906 4140
rect 272426 4128 272432 4140
rect 253900 4100 272432 4128
rect 253900 4088 253906 4100
rect 272426 4088 272432 4100
rect 272484 4088 272490 4140
rect 329190 4088 329196 4140
rect 329248 4128 329254 4140
rect 347222 4128 347228 4140
rect 329248 4100 347228 4128
rect 329248 4088 329254 4100
rect 347222 4088 347228 4100
rect 347280 4088 347286 4140
rect 249702 4020 249708 4072
rect 249760 4060 249766 4072
rect 268838 4060 268844 4072
rect 249760 4032 268844 4060
rect 249760 4020 249766 4032
rect 268838 4020 268844 4032
rect 268896 4020 268902 4072
rect 327994 4020 328000 4072
rect 328052 4060 328058 4072
rect 346670 4060 346676 4072
rect 328052 4032 346676 4060
rect 328052 4020 328058 4032
rect 346670 4020 346676 4032
rect 346728 4020 346734 4072
rect 259178 3952 259184 4004
rect 259236 3992 259242 4004
rect 281902 3992 281908 4004
rect 259236 3964 281908 3992
rect 259236 3952 259242 3964
rect 281902 3952 281908 3964
rect 281960 3952 281966 4004
rect 325602 3952 325608 4004
rect 325660 3992 325666 4004
rect 344370 3992 344376 4004
rect 325660 3964 344376 3992
rect 325660 3952 325666 3964
rect 344370 3952 344376 3964
rect 344428 3952 344434 4004
rect 128170 3884 128176 3936
rect 128228 3924 128234 3936
rect 182910 3924 182916 3936
rect 128228 3896 182916 3924
rect 128228 3884 128234 3896
rect 182910 3884 182916 3896
rect 182968 3884 182974 3936
rect 251082 3884 251088 3936
rect 251140 3924 251146 3936
rect 276014 3924 276020 3936
rect 251140 3896 276020 3924
rect 251140 3884 251146 3896
rect 276014 3884 276020 3896
rect 276072 3884 276078 3936
rect 324406 3884 324412 3936
rect 324464 3924 324470 3936
rect 346762 3924 346768 3936
rect 324464 3896 346768 3924
rect 324464 3884 324470 3896
rect 346762 3884 346768 3896
rect 346820 3884 346826 3936
rect 141234 3816 141240 3868
rect 141292 3856 141298 3868
rect 197354 3856 197360 3868
rect 141292 3828 197360 3856
rect 141292 3816 141298 3828
rect 197354 3816 197360 3828
rect 197412 3816 197418 3868
rect 203886 3816 203892 3868
rect 203944 3856 203950 3868
rect 243538 3856 243544 3868
rect 203944 3828 243544 3856
rect 203944 3816 203950 3828
rect 243538 3816 243544 3828
rect 243596 3816 243602 3868
rect 257614 3816 257620 3868
rect 257672 3856 257678 3868
rect 285398 3856 285404 3868
rect 257672 3828 285404 3856
rect 257672 3816 257678 3828
rect 285398 3816 285404 3828
rect 285456 3816 285462 3868
rect 322106 3816 322112 3868
rect 322164 3856 322170 3868
rect 345842 3856 345848 3868
rect 322164 3828 345848 3856
rect 322164 3816 322170 3828
rect 345842 3816 345848 3828
rect 345900 3816 345906 3868
rect 70302 3748 70308 3800
rect 70360 3788 70366 3800
rect 127618 3788 127624 3800
rect 70360 3760 127624 3788
rect 70360 3748 70366 3760
rect 127618 3748 127624 3760
rect 127676 3748 127682 3800
rect 175458 3748 175464 3800
rect 175516 3788 175522 3800
rect 249058 3788 249064 3800
rect 175516 3760 249064 3788
rect 175516 3748 175522 3760
rect 249058 3748 249064 3760
rect 249116 3748 249122 3800
rect 257706 3748 257712 3800
rect 257764 3788 257770 3800
rect 288986 3788 288992 3800
rect 257764 3760 288992 3788
rect 257764 3748 257770 3760
rect 288986 3748 288992 3760
rect 289044 3748 289050 3800
rect 320910 3748 320916 3800
rect 320968 3788 320974 3800
rect 343910 3788 343916 3800
rect 320968 3760 343916 3788
rect 320968 3748 320974 3760
rect 343910 3748 343916 3760
rect 343968 3748 343974 3800
rect 86862 3680 86868 3732
rect 86920 3720 86926 3732
rect 181438 3720 181444 3732
rect 86920 3692 181444 3720
rect 86920 3680 86926 3692
rect 181438 3680 181444 3692
rect 181496 3680 181502 3732
rect 196802 3680 196808 3732
rect 196860 3720 196866 3732
rect 243630 3720 243636 3732
rect 196860 3692 243636 3720
rect 196860 3680 196866 3692
rect 243630 3680 243636 3692
rect 243688 3680 243694 3732
rect 244182 3680 244188 3732
rect 244240 3720 244246 3732
rect 278314 3720 278320 3732
rect 244240 3692 278320 3720
rect 244240 3680 244246 3692
rect 278314 3680 278320 3692
rect 278372 3680 278378 3732
rect 326798 3680 326804 3732
rect 326856 3720 326862 3732
rect 349522 3720 349528 3732
rect 326856 3692 349528 3720
rect 326856 3680 326862 3692
rect 349522 3680 349528 3692
rect 349580 3680 349586 3732
rect 65518 3612 65524 3664
rect 65576 3652 65582 3664
rect 196066 3652 196072 3664
rect 65576 3624 196072 3652
rect 65576 3612 65582 3624
rect 196066 3612 196072 3624
rect 196124 3612 196130 3664
rect 200298 3612 200304 3664
rect 200356 3652 200362 3664
rect 242158 3652 242164 3664
rect 200356 3624 242164 3652
rect 200356 3612 200362 3624
rect 242158 3612 242164 3624
rect 242216 3612 242222 3664
rect 259362 3612 259368 3664
rect 259420 3652 259426 3664
rect 296070 3652 296076 3664
rect 259420 3624 296076 3652
rect 259420 3612 259426 3624
rect 296070 3612 296076 3624
rect 296128 3612 296134 3664
rect 323302 3612 323308 3664
rect 323360 3652 323366 3664
rect 348142 3652 348148 3664
rect 323360 3624 348148 3652
rect 323360 3612 323366 3624
rect 348142 3612 348148 3624
rect 348200 3612 348206 3664
rect 2866 3544 2872 3596
rect 2924 3584 2930 3596
rect 175918 3584 175924 3596
rect 2924 3556 175924 3584
rect 2924 3544 2930 3556
rect 175918 3544 175924 3556
rect 175976 3544 175982 3596
rect 179046 3544 179052 3596
rect 179104 3584 179110 3596
rect 233878 3584 233884 3596
rect 179104 3556 233884 3584
rect 179104 3544 179110 3556
rect 233878 3544 233884 3556
rect 233936 3544 233942 3596
rect 244918 3544 244924 3596
rect 244976 3544 244982 3596
rect 256602 3544 256608 3596
rect 256660 3584 256666 3596
rect 292574 3584 292580 3596
rect 256660 3556 292580 3584
rect 256660 3544 256666 3556
rect 292574 3544 292580 3556
rect 292632 3544 292638 3596
rect 318518 3544 318524 3596
rect 318576 3584 318582 3596
rect 344646 3584 344652 3596
rect 318576 3556 344652 3584
rect 318576 3544 318582 3556
rect 344646 3544 344652 3556
rect 344704 3544 344710 3596
rect 349614 3584 349620 3596
rect 344986 3556 349620 3584
rect 30098 3476 30104 3528
rect 30156 3516 30162 3528
rect 221458 3516 221464 3528
rect 30156 3488 221464 3516
rect 30156 3476 30162 3488
rect 221458 3476 221464 3488
rect 221516 3476 221522 3528
rect 226334 3476 226340 3528
rect 226392 3516 226398 3528
rect 227530 3516 227536 3528
rect 226392 3488 227536 3516
rect 226392 3476 226398 3488
rect 227530 3476 227536 3488
rect 227588 3476 227594 3528
rect 227622 3476 227628 3528
rect 227680 3516 227686 3528
rect 242250 3516 242256 3528
rect 227680 3488 242256 3516
rect 227680 3476 227686 3488
rect 242250 3476 242256 3488
rect 242308 3476 242314 3528
rect 15930 3408 15936 3460
rect 15988 3448 15994 3460
rect 244936 3448 244964 3544
rect 254670 3476 254676 3528
rect 254728 3516 254734 3528
rect 256050 3516 256056 3528
rect 254728 3488 256056 3516
rect 254728 3476 254734 3488
rect 256050 3476 256056 3488
rect 256108 3476 256114 3528
rect 257522 3476 257528 3528
rect 257580 3516 257586 3528
rect 299658 3516 299664 3528
rect 257580 3488 299664 3516
rect 257580 3476 257586 3488
rect 299658 3476 299664 3488
rect 299716 3476 299722 3528
rect 319714 3476 319720 3528
rect 319772 3516 319778 3528
rect 344986 3516 345014 3556
rect 349614 3544 349620 3556
rect 349672 3544 349678 3596
rect 319772 3488 345014 3516
rect 319772 3476 319778 3488
rect 365806 3476 365812 3528
rect 365864 3516 365870 3528
rect 367002 3516 367008 3528
rect 365864 3488 367008 3516
rect 365864 3476 365870 3488
rect 367002 3476 367008 3488
rect 367060 3476 367066 3528
rect 374086 3476 374092 3528
rect 374144 3516 374150 3528
rect 375282 3516 375288 3528
rect 374144 3488 375288 3516
rect 374144 3476 374150 3488
rect 375282 3476 375288 3488
rect 375340 3476 375346 3528
rect 382366 3476 382372 3528
rect 382424 3516 382430 3528
rect 383562 3516 383568 3528
rect 382424 3488 383568 3516
rect 382424 3476 382430 3488
rect 383562 3476 383568 3488
rect 383620 3476 383626 3528
rect 390646 3476 390652 3528
rect 390704 3516 390710 3528
rect 391842 3516 391848 3528
rect 390704 3488 391848 3516
rect 390704 3476 390710 3488
rect 391842 3476 391848 3488
rect 391900 3476 391906 3528
rect 407206 3476 407212 3528
rect 407264 3516 407270 3528
rect 408402 3516 408408 3528
rect 407264 3488 408408 3516
rect 407264 3476 407270 3488
rect 408402 3476 408408 3488
rect 408460 3476 408466 3528
rect 415486 3476 415492 3528
rect 415544 3516 415550 3528
rect 416682 3516 416688 3528
rect 415544 3488 416688 3516
rect 415544 3476 415550 3488
rect 416682 3476 416688 3488
rect 416740 3476 416746 3528
rect 423766 3476 423772 3528
rect 423824 3516 423830 3528
rect 424962 3516 424968 3528
rect 423824 3488 424968 3516
rect 423824 3476 423830 3488
rect 424962 3476 424968 3488
rect 425020 3476 425026 3528
rect 432046 3476 432052 3528
rect 432104 3516 432110 3528
rect 433242 3516 433248 3528
rect 432104 3488 433248 3516
rect 432104 3476 432110 3488
rect 433242 3476 433248 3488
rect 433300 3476 433306 3528
rect 448606 3476 448612 3528
rect 448664 3516 448670 3528
rect 449802 3516 449808 3528
rect 448664 3488 449808 3516
rect 448664 3476 448670 3488
rect 449802 3476 449808 3488
rect 449860 3476 449866 3528
rect 456886 3476 456892 3528
rect 456944 3516 456950 3528
rect 458082 3516 458088 3528
rect 456944 3488 458088 3516
rect 456944 3476 456950 3488
rect 458082 3476 458088 3488
rect 458140 3476 458146 3528
rect 465074 3476 465080 3528
rect 465132 3516 465138 3528
rect 465902 3516 465908 3528
rect 465132 3488 465908 3516
rect 465132 3476 465138 3488
rect 465902 3476 465908 3488
rect 465960 3476 465966 3528
rect 489914 3476 489920 3528
rect 489972 3516 489978 3528
rect 490742 3516 490748 3528
rect 489972 3488 490748 3516
rect 489972 3476 489978 3488
rect 490742 3476 490748 3488
rect 490800 3476 490806 3528
rect 498194 3476 498200 3528
rect 498252 3516 498258 3528
rect 499022 3516 499028 3528
rect 498252 3488 499028 3516
rect 498252 3476 498258 3488
rect 499022 3476 499028 3488
rect 499080 3476 499086 3528
rect 514754 3476 514760 3528
rect 514812 3516 514818 3528
rect 515582 3516 515588 3528
rect 514812 3488 515588 3516
rect 514812 3476 514818 3488
rect 515582 3476 515588 3488
rect 515640 3476 515646 3528
rect 523034 3476 523040 3528
rect 523092 3516 523098 3528
rect 523862 3516 523868 3528
rect 523092 3488 523868 3516
rect 523092 3476 523098 3488
rect 523862 3476 523868 3488
rect 523920 3476 523926 3528
rect 539594 3476 539600 3528
rect 539652 3516 539658 3528
rect 540422 3516 540428 3528
rect 539652 3488 540428 3516
rect 539652 3476 539658 3488
rect 540422 3476 540428 3488
rect 540480 3476 540486 3528
rect 547874 3476 547880 3528
rect 547932 3516 547938 3528
rect 548702 3516 548708 3528
rect 547932 3488 548708 3516
rect 547932 3476 547938 3488
rect 548702 3476 548708 3488
rect 548760 3476 548766 3528
rect 580994 3476 581000 3528
rect 581052 3516 581058 3528
rect 581822 3516 581828 3528
rect 581052 3488 581828 3516
rect 581052 3476 581058 3488
rect 581822 3476 581828 3488
rect 581880 3476 581886 3528
rect 15988 3420 244964 3448
rect 15988 3408 15994 3420
rect 246390 3408 246396 3460
rect 246448 3448 246454 3460
rect 254578 3448 254584 3460
rect 246448 3420 254584 3448
rect 246448 3408 246454 3420
rect 254578 3408 254584 3420
rect 254636 3408 254642 3460
rect 257430 3408 257436 3460
rect 257488 3448 257494 3460
rect 303154 3448 303160 3460
rect 257488 3420 303160 3448
rect 257488 3408 257494 3420
rect 303154 3408 303160 3420
rect 303212 3408 303218 3460
rect 315022 3408 315028 3460
rect 315080 3448 315086 3460
rect 346394 3448 346400 3460
rect 315080 3420 346400 3448
rect 315080 3408 315086 3420
rect 346394 3408 346400 3420
rect 346452 3408 346458 3460
rect 356698 3408 356704 3460
rect 356756 3448 356762 3460
rect 579798 3448 579804 3460
rect 356756 3420 579804 3448
rect 356756 3408 356762 3420
rect 579798 3408 579804 3420
rect 579856 3408 579862 3460
rect 44174 3340 44180 3392
rect 44232 3380 44238 3392
rect 45094 3380 45100 3392
rect 44232 3352 45100 3380
rect 44232 3340 44238 3352
rect 45094 3340 45100 3352
rect 45152 3340 45158 3392
rect 259086 3340 259092 3392
rect 259144 3380 259150 3392
rect 271230 3380 271236 3392
rect 259144 3352 271236 3380
rect 259144 3340 259150 3352
rect 271230 3340 271236 3352
rect 271288 3340 271294 3392
rect 330386 3340 330392 3392
rect 330444 3380 330450 3392
rect 347866 3380 347872 3392
rect 330444 3352 347872 3380
rect 330444 3340 330450 3352
rect 347866 3340 347872 3352
rect 347924 3340 347930 3392
rect 253750 3272 253756 3324
rect 253808 3312 253814 3324
rect 265342 3312 265348 3324
rect 253808 3284 265348 3312
rect 253808 3272 253814 3284
rect 265342 3272 265348 3284
rect 265400 3272 265406 3324
rect 331582 3272 331588 3324
rect 331640 3312 331646 3324
rect 346578 3312 346584 3324
rect 331640 3284 346584 3312
rect 331640 3272 331646 3284
rect 346578 3272 346584 3284
rect 346636 3272 346642 3324
rect 259270 3204 259276 3256
rect 259328 3244 259334 3256
rect 267734 3244 267740 3256
rect 259328 3216 267740 3244
rect 259328 3204 259334 3216
rect 267734 3204 267740 3216
rect 267792 3204 267798 3256
rect 332686 3204 332692 3256
rect 332744 3244 332750 3256
rect 346854 3244 346860 3256
rect 332744 3216 346860 3244
rect 332744 3204 332750 3216
rect 346854 3204 346860 3216
rect 346912 3204 346918 3256
rect 252370 3136 252376 3188
rect 252428 3176 252434 3188
rect 255958 3176 255964 3188
rect 252428 3148 255964 3176
rect 252428 3136 252434 3148
rect 255958 3136 255964 3148
rect 256016 3136 256022 3188
rect 226334 2796 226340 2848
rect 226392 2836 226398 2848
rect 227622 2836 227628 2848
rect 226392 2808 227628 2836
rect 226392 2796 226398 2808
rect 227622 2796 227628 2808
rect 227680 2796 227686 2848
rect 357434 2184 357440 2236
rect 357492 2224 357498 2236
rect 358722 2224 358728 2236
rect 357492 2196 358728 2224
rect 357492 2184 357498 2196
rect 358722 2184 358728 2196
rect 358780 2184 358786 2236
rect 398834 2184 398840 2236
rect 398892 2224 398898 2236
rect 400122 2224 400128 2236
rect 398892 2196 400128 2224
rect 398892 2184 398898 2196
rect 400122 2184 400128 2196
rect 400180 2184 400186 2236
rect 440234 2184 440240 2236
rect 440292 2224 440298 2236
rect 441522 2224 441528 2236
rect 440292 2196 441528 2224
rect 440292 2184 440298 2196
rect 441522 2184 441528 2196
rect 441580 2184 441586 2236
<< via1 >>
rect 71780 702992 71832 703044
rect 72976 702992 73028 703044
rect 201500 702992 201552 703044
rect 202788 702992 202840 703044
rect 170312 700476 170364 700528
rect 192484 700476 192536 700528
rect 255596 700476 255648 700528
rect 283840 700476 283892 700528
rect 331864 700476 331916 700528
rect 397460 700476 397512 700528
rect 154120 700408 154172 700460
rect 242164 700408 242216 700460
rect 265624 700408 265676 700460
rect 348792 700408 348844 700460
rect 89168 700340 89220 700392
rect 257620 700340 257672 700392
rect 324964 700340 325016 700392
rect 332508 700340 332560 700392
rect 347044 700340 347096 700392
rect 462320 700340 462372 700392
rect 24308 700272 24360 700324
rect 192576 700272 192628 700324
rect 258724 700272 258776 700324
rect 413652 700272 413704 700324
rect 218980 699660 219032 699712
rect 220084 699660 220136 699712
rect 266360 697552 266412 697604
rect 267648 697552 267700 697604
rect 264244 696940 264296 696992
rect 580172 696940 580224 696992
rect 3424 683204 3476 683256
rect 257344 683204 257396 683256
rect 253204 683136 253256 683188
rect 580172 683136 580224 683188
rect 3424 670760 3476 670812
rect 258816 670760 258868 670812
rect 251824 670692 251876 670744
rect 580172 670692 580224 670744
rect 3424 656888 3476 656940
rect 192668 656888 192720 656940
rect 261484 643084 261536 643136
rect 580172 643084 580224 643136
rect 3424 632068 3476 632120
rect 259828 632068 259880 632120
rect 249892 630640 249944 630692
rect 580172 630640 580224 630692
rect 2780 619080 2832 619132
rect 4804 619080 4856 619132
rect 251916 616836 251968 616888
rect 580172 616836 580224 616888
rect 3240 605820 3292 605872
rect 259552 605820 259604 605872
rect 261576 590656 261628 590708
rect 579804 590656 579856 590708
rect 136640 590044 136692 590096
rect 256792 590044 256844 590096
rect 104900 589976 104952 590028
rect 257436 589976 257488 590028
rect 252652 589908 252704 589960
rect 429200 589908 429252 589960
rect 2780 566040 2832 566092
rect 4896 566040 4948 566092
rect 2780 553664 2832 553716
rect 4988 553664 5040 553716
rect 279424 536800 279476 536852
rect 376944 536800 376996 536852
rect 278044 535440 278096 535492
rect 377036 535440 377088 535492
rect 278136 534080 278188 534132
rect 376944 534080 376996 534132
rect 275284 532720 275336 532772
rect 377036 532720 377088 532772
rect 278228 531292 278280 531344
rect 376944 531292 376996 531344
rect 273904 529932 273956 529984
rect 376944 529932 376996 529984
rect 273996 528572 274048 528624
rect 376852 528572 376904 528624
rect 471244 510620 471296 510672
rect 579620 510620 579672 510672
rect 295984 509260 296036 509312
rect 376944 509260 376996 509312
rect 296076 507900 296128 507952
rect 376760 507900 376812 507952
rect 271144 507832 271196 507884
rect 377036 507832 377088 507884
rect 3332 501304 3384 501356
rect 7564 501304 7616 501356
rect 123392 498040 123444 498092
rect 124864 498040 124916 498092
rect 287428 497156 287480 497208
rect 397460 497156 397512 497208
rect 288624 497088 288676 497140
rect 398840 497088 398892 497140
rect 119344 497020 119396 497072
rect 279700 497020 279752 497072
rect 288532 497020 288584 497072
rect 398932 497020 398984 497072
rect 126796 496952 126848 497004
rect 282184 496952 282236 497004
rect 292672 496952 292724 497004
rect 403164 496952 403216 497004
rect 125232 496884 125284 496936
rect 285220 496884 285272 496936
rect 285772 496884 285824 496936
rect 404360 496884 404412 496936
rect 115480 496816 115532 496868
rect 116584 496816 116636 496868
rect 287152 496816 287204 496868
rect 409880 496816 409932 496868
rect 249156 484372 249208 484424
rect 580172 484372 580224 484424
rect 3332 474716 3384 474768
rect 261668 474716 261720 474768
rect 247132 470568 247184 470620
rect 579988 470568 580040 470620
rect 3332 462340 3384 462392
rect 175924 462340 175976 462392
rect 247408 456764 247460 456816
rect 580172 456764 580224 456816
rect 3332 448536 3384 448588
rect 262588 448536 262640 448588
rect 245752 430584 245804 430636
rect 579620 430584 579672 430636
rect 97540 426368 97592 426420
rect 295616 426368 295668 426420
rect 296076 426368 296128 426420
rect 3148 422288 3200 422340
rect 261760 422288 261812 422340
rect 247224 418140 247276 418192
rect 579712 418140 579764 418192
rect 155868 414808 155920 414860
rect 284392 414808 284444 414860
rect 151728 414740 151780 414792
rect 283656 414740 283708 414792
rect 146208 414672 146260 414724
rect 281908 414672 281960 414724
rect 291292 414672 291344 414724
rect 401600 414672 401652 414724
rect 3148 409844 3200 409896
rect 234528 409844 234580 409896
rect 263784 409844 263836 409896
rect 248512 406376 248564 406428
rect 580356 406376 580408 406428
rect 246028 404336 246080 404388
rect 579988 404336 580040 404388
rect 124864 401004 124916 401056
rect 283012 401004 283064 401056
rect 121276 400936 121328 400988
rect 281816 400936 281868 400988
rect 122748 400868 122800 400920
rect 283104 400868 283156 400920
rect 254032 399712 254084 399764
rect 266360 399712 266412 399764
rect 161388 399644 161440 399696
rect 285864 399644 285916 399696
rect 140688 399576 140740 399628
rect 280252 399576 280304 399628
rect 118608 399508 118660 399560
rect 278596 399508 278648 399560
rect 121368 399440 121420 399492
rect 280804 399440 280856 399492
rect 136548 398148 136600 398200
rect 280344 398148 280396 398200
rect 97816 398080 97868 398132
rect 277308 398080 277360 398132
rect 3332 397468 3384 397520
rect 263416 397468 263468 397520
rect 97632 397400 97684 397452
rect 295984 397400 296036 397452
rect 99104 397332 99156 397384
rect 275284 397332 275336 397384
rect 131028 396788 131080 396840
rect 279148 396788 279200 396840
rect 99196 396720 99248 396772
rect 275928 396720 275980 396772
rect 294052 396720 294104 396772
rect 405740 396720 405792 396772
rect 275376 396040 275428 396092
rect 275928 396040 275980 396092
rect 278136 396040 278188 396092
rect 98920 395972 98972 396024
rect 273996 395972 274048 396024
rect 99012 395904 99064 395956
rect 273904 395904 273956 395956
rect 274180 395904 274232 395956
rect 277308 395904 277360 395956
rect 279424 395904 279476 395956
rect 294144 395428 294196 395480
rect 404452 395428 404504 395480
rect 116584 395360 116636 395412
rect 271972 395360 272024 395412
rect 290740 395360 290792 395412
rect 400220 395360 400272 395412
rect 114468 395292 114520 395344
rect 272524 395292 272576 395344
rect 294604 395292 294656 395344
rect 440240 395292 440292 395344
rect 254584 394136 254636 394188
rect 265624 394136 265676 394188
rect 242164 394068 242216 394120
rect 257160 394068 257212 394120
rect 291384 394068 291436 394120
rect 425060 394068 425112 394120
rect 113088 394000 113140 394052
rect 272616 394000 272668 394052
rect 292396 394000 292448 394052
rect 429200 394000 429252 394052
rect 3608 393932 3660 393984
rect 262128 393932 262180 393984
rect 293500 393932 293552 393984
rect 434720 393932 434772 393984
rect 233792 393320 233844 393372
rect 260472 393388 260524 393440
rect 252928 393320 252980 393372
rect 258724 393320 258776 393372
rect 220084 392844 220136 392896
rect 256240 392844 256292 392896
rect 253020 392776 253072 392828
rect 477500 392776 477552 392828
rect 7564 392708 7616 392760
rect 261944 392708 261996 392760
rect 251272 392640 251324 392692
rect 542360 392640 542412 392692
rect 192576 392572 192628 392624
rect 233976 392572 234028 392624
rect 248788 392572 248840 392624
rect 580540 392572 580592 392624
rect 248512 392436 248564 392488
rect 249616 392436 249668 392488
rect 233976 391960 234028 392012
rect 258724 391960 258776 392012
rect 192668 391552 192720 391604
rect 259276 391552 259328 391604
rect 254400 391484 254452 391536
rect 324964 391484 325016 391536
rect 253480 391416 253532 391468
rect 331864 391416 331916 391468
rect 252744 391348 252796 391400
rect 347044 391348 347096 391400
rect 6920 391280 6972 391332
rect 258540 391280 258592 391332
rect 4988 391212 5040 391264
rect 260932 391212 260984 391264
rect 251364 390532 251416 390584
rect 253204 390532 253256 390584
rect 258816 390532 258868 390584
rect 260196 390532 260248 390584
rect 273076 390464 273128 390516
rect 394700 390464 394752 390516
rect 250168 390124 250220 390176
rect 261484 390124 261536 390176
rect 249340 390056 249392 390108
rect 261576 390056 261628 390108
rect 250996 389988 251048 390040
rect 264244 389988 264296 390040
rect 271972 389988 272024 390040
rect 273076 389988 273128 390040
rect 71780 389920 71832 389972
rect 257620 389920 257672 389972
rect 252008 389852 252060 389904
rect 527180 389852 527232 389904
rect 248420 389784 248472 389836
rect 580448 389784 580500 389836
rect 287152 389716 287204 389768
rect 287980 389716 288032 389768
rect 288532 389308 288584 389360
rect 289636 389308 289688 389360
rect 254952 388832 255004 388884
rect 299480 388832 299532 388884
rect 201500 388764 201552 388816
rect 255964 388764 256016 388816
rect 254308 388696 254360 388748
rect 364340 388696 364392 388748
rect 40040 388628 40092 388680
rect 258172 388628 258224 388680
rect 252468 388560 252520 388612
rect 494060 388560 494112 388612
rect 4896 388492 4948 388544
rect 261300 388492 261352 388544
rect 3516 388424 3568 388476
rect 261484 388424 261536 388476
rect 283012 388424 283064 388476
rect 284116 388424 284168 388476
rect 285772 388424 285824 388476
rect 286876 388424 286928 388476
rect 294052 388424 294104 388476
rect 295156 388424 295208 388476
rect 290188 388356 290240 388408
rect 419540 388424 419592 388476
rect 234620 387404 234672 387456
rect 255688 387404 255740 387456
rect 192484 387336 192536 387388
rect 256516 387336 256568 387388
rect 248328 387268 248380 387320
rect 471244 387268 471296 387320
rect 3424 387200 3476 387252
rect 260656 387200 260708 387252
rect 251640 387132 251692 387184
rect 558920 387132 558972 387184
rect 249248 387064 249300 387116
rect 580264 387064 580316 387116
rect 249984 386520 250036 386572
rect 251916 386520 251968 386572
rect 261760 386520 261812 386572
rect 263140 386520 263192 386572
rect 247776 386452 247828 386504
rect 249156 386452 249208 386504
rect 250812 386452 250864 386504
rect 251824 386452 251876 386504
rect 257344 386452 257396 386504
rect 259000 386452 259052 386504
rect 261668 386452 261720 386504
rect 262312 386452 262364 386504
rect 235816 386384 235868 386436
rect 281632 386452 281684 386504
rect 275376 386384 275428 386436
rect 275836 386384 275888 386436
rect 97724 386316 97776 386368
rect 271512 386316 271564 386368
rect 272524 386248 272576 386300
rect 272800 386248 272852 386300
rect 393320 386316 393372 386368
rect 272248 386180 272300 386232
rect 272616 386180 272668 386232
rect 391940 386248 391992 386300
rect 175924 385840 175976 385892
rect 235540 385840 235592 385892
rect 125508 385772 125560 385824
rect 278136 385772 278188 385824
rect 99288 385704 99340 385756
rect 274824 385704 274876 385756
rect 278228 385704 278280 385756
rect 97908 385636 97960 385688
rect 276480 385636 276532 385688
rect 278044 385636 278096 385688
rect 289268 385636 289320 385688
rect 415400 385636 415452 385688
rect 244924 385296 244976 385348
rect 253848 385296 253900 385348
rect 247132 385228 247184 385280
rect 247960 385228 248012 385280
rect 251272 385228 251324 385280
rect 252100 385228 252152 385280
rect 252652 385228 252704 385280
rect 253204 385228 253256 385280
rect 235540 385160 235592 385212
rect 235724 385160 235776 385212
rect 262864 385228 262916 385280
rect 254032 385160 254084 385212
rect 255136 385160 255188 385212
rect 259552 385160 259604 385212
rect 260104 385160 260156 385212
rect 280252 385160 280304 385212
rect 281356 385160 281408 385212
rect 252928 385092 252980 385144
rect 253756 385092 253808 385144
rect 253848 385092 253900 385144
rect 577964 385092 578016 385144
rect 244096 385024 244148 385076
rect 577780 385024 577832 385076
rect 282184 384956 282236 385008
rect 286324 384956 286376 385008
rect 241060 384820 241112 384872
rect 295340 384820 295392 384872
rect 236828 384752 236880 384804
rect 267004 384752 267056 384804
rect 286784 384752 286836 384804
rect 296812 384752 296864 384804
rect 246396 384684 246448 384736
rect 293776 384684 293828 384736
rect 174544 384616 174596 384668
rect 270316 384616 270368 384668
rect 285588 384616 285640 384668
rect 301872 384616 301924 384668
rect 243820 384548 243872 384600
rect 579988 384548 580040 384600
rect 242808 384480 242860 384532
rect 580540 384480 580592 384532
rect 267648 384412 267700 384464
rect 291844 384412 291896 384464
rect 235632 384344 235684 384396
rect 269764 384344 269816 384396
rect 264888 384276 264940 384328
rect 301780 384276 301832 384328
rect 231124 384208 231176 384260
rect 269488 384208 269540 384260
rect 279516 384208 279568 384260
rect 344652 384208 344704 384260
rect 274456 384140 274508 384192
rect 300124 384140 300176 384192
rect 241336 384072 241388 384124
rect 289728 384072 289780 384124
rect 291292 384072 291344 384124
rect 291844 384072 291896 384124
rect 240048 384004 240100 384056
rect 290924 384004 290976 384056
rect 291752 384004 291804 384056
rect 300492 384072 300544 384124
rect 296536 384004 296588 384056
rect 344284 384004 344336 384056
rect 233976 383936 234028 383988
rect 275560 383936 275612 383988
rect 293408 383936 293460 383988
rect 344100 383936 344152 383988
rect 248880 383868 248932 383920
rect 264520 383868 264572 383920
rect 285128 383868 285180 383920
rect 347780 383868 347832 383920
rect 245200 383800 245252 383852
rect 261208 383800 261260 383852
rect 290648 383800 290700 383852
rect 300216 383800 300268 383852
rect 239404 383732 239456 383784
rect 270040 383732 270092 383784
rect 292764 383732 292816 383784
rect 301504 383732 301556 383784
rect 261300 383664 261352 383716
rect 274548 383664 274600 383716
rect 283564 383664 283616 383716
rect 291108 383664 291160 383716
rect 294512 383664 294564 383716
rect 300400 383664 300452 383716
rect 245660 383256 245712 383308
rect 248880 383256 248932 383308
rect 244648 383188 244700 383240
rect 245476 383120 245528 383172
rect 249064 383188 249116 383240
rect 577596 383188 577648 383240
rect 235448 383052 235500 383104
rect 578056 383120 578108 383172
rect 580264 383052 580316 383104
rect 264796 382984 264848 383036
rect 3792 382916 3844 382968
rect 245660 382916 245712 382968
rect 245752 382916 245804 382968
rect 246856 382916 246908 382968
rect 258632 382916 258684 382968
rect 264060 382916 264112 382968
rect 264888 382916 264940 382968
rect 291108 382916 291160 382968
rect 322940 382916 322992 382968
rect 235172 382848 235224 382900
rect 264244 382848 264296 382900
rect 234160 382780 234212 382832
rect 275008 382780 275060 382832
rect 278964 382780 279016 382832
rect 301688 382780 301740 382832
rect 234252 382712 234304 382764
rect 280528 382712 280580 382764
rect 246120 382644 246172 382696
rect 300768 382644 300820 382696
rect 174636 382576 174688 382628
rect 258632 382576 258684 382628
rect 284484 382576 284536 382628
rect 337384 382576 337436 382628
rect 94504 382508 94556 382560
rect 267832 382508 267884 382560
rect 286140 382508 286192 382560
rect 349252 382508 349304 382560
rect 91744 382440 91796 382492
rect 266176 382440 266228 382492
rect 272524 382440 272576 382492
rect 347872 382440 347924 382492
rect 233792 382372 233844 382424
rect 265348 382372 265400 382424
rect 289084 382372 289136 382424
rect 301596 382372 301648 382424
rect 235356 382304 235408 382356
rect 265072 382304 265124 382356
rect 287244 382304 287296 382356
rect 300308 382304 300360 382356
rect 232504 382236 232556 382288
rect 265624 382236 265676 382288
rect 280068 382236 280120 382288
rect 299480 382236 299532 382288
rect 242992 381896 243044 381948
rect 248236 381896 248288 381948
rect 241612 381828 241664 381880
rect 257068 381964 257120 382016
rect 263968 381964 264020 382016
rect 265900 381964 265952 382016
rect 252928 381896 252980 381948
rect 267280 381896 267332 381948
rect 245752 381760 245804 381812
rect 256240 381760 256292 381812
rect 3700 381556 3752 381608
rect 236828 381692 236880 381744
rect 243544 381692 243596 381744
rect 247408 381692 247460 381744
rect 247684 381692 247736 381744
rect 250720 381692 250772 381744
rect 255136 381692 255188 381744
rect 259828 381692 259880 381744
rect 235908 381624 235960 381676
rect 235540 381556 235592 381608
rect 252928 381556 252980 381608
rect 3424 381488 3476 381540
rect 239404 381488 239456 381540
rect 234436 381216 234488 381268
rect 247684 381488 247736 381540
rect 250720 381488 250772 381540
rect 268936 381828 268988 381880
rect 261208 381624 261260 381676
rect 270592 381692 270644 381744
rect 241612 381420 241664 381472
rect 242992 381420 243044 381472
rect 244372 381420 244424 381472
rect 247408 381420 247460 381472
rect 90456 381080 90508 381132
rect 3608 381012 3660 381064
rect 248236 381420 248288 381472
rect 255136 381420 255188 381472
rect 256240 381420 256292 381472
rect 257068 381420 257120 381472
rect 259828 381420 259880 381472
rect 276940 381624 276992 381676
rect 282184 381624 282236 381676
rect 263968 381420 264020 381472
rect 266728 381420 266780 381472
rect 271972 381420 272024 381472
rect 277492 381488 277544 381540
rect 296812 381624 296864 381676
rect 306380 381624 306432 381676
rect 293776 381556 293828 381608
rect 579896 381556 579948 381608
rect 276940 381420 276992 381472
rect 580080 381488 580132 381540
rect 282184 381420 282236 381472
rect 283012 381420 283064 381472
rect 300952 381216 301004 381268
rect 301964 381148 302016 381200
rect 300860 381080 300912 381132
rect 344008 381012 344060 381064
rect 580724 380944 580776 380996
rect 580908 380876 580960 380928
rect 300768 379448 300820 379500
rect 580172 379448 580224 379500
rect 579988 378768 580040 378820
rect 580816 378768 580868 378820
rect 3148 372512 3200 372564
rect 174636 372512 174688 372564
rect 301964 353200 302016 353252
rect 579988 353200 580040 353252
rect 2964 346332 3016 346384
rect 235172 346332 235224 346384
rect 244096 338512 244148 338564
rect 244740 338036 244792 338088
rect 242992 337968 243044 338020
rect 244464 337900 244516 337952
rect 245614 337900 245666 337952
rect 245706 337900 245758 337952
rect 245890 337900 245942 337952
rect 246258 337900 246310 337952
rect 246442 337900 246494 337952
rect 246718 337900 246770 337952
rect 246810 337900 246862 337952
rect 246902 337900 246954 337952
rect 247086 337900 247138 337952
rect 247178 337900 247230 337952
rect 247362 337900 247414 337952
rect 245108 337832 245160 337884
rect 244280 337764 244332 337816
rect 245522 337764 245574 337816
rect 245936 337696 245988 337748
rect 246028 337628 246080 337680
rect 246626 337832 246678 337884
rect 246672 337696 246724 337748
rect 246764 337696 246816 337748
rect 246580 337560 246632 337612
rect 246488 337492 246540 337544
rect 245016 337424 245068 337476
rect 247270 337832 247322 337884
rect 247822 337900 247874 337952
rect 247132 337764 247184 337816
rect 247638 337832 247690 337884
rect 247408 337764 247460 337816
rect 248282 337900 248334 337952
rect 248374 337900 248426 337952
rect 248650 337900 248702 337952
rect 248742 337900 248794 337952
rect 248834 337900 248886 337952
rect 248926 337900 248978 337952
rect 249110 337900 249162 337952
rect 249202 337900 249254 337952
rect 249294 337900 249346 337952
rect 248006 337832 248058 337884
rect 248098 337832 248150 337884
rect 247224 337696 247276 337748
rect 247316 337696 247368 337748
rect 247224 337560 247276 337612
rect 247868 337764 247920 337816
rect 247592 337628 247644 337680
rect 247776 337560 247828 337612
rect 248466 337832 248518 337884
rect 248512 337696 248564 337748
rect 248788 337764 248840 337816
rect 248880 337696 248932 337748
rect 248328 337628 248380 337680
rect 248604 337628 248656 337680
rect 249156 337628 249208 337680
rect 249248 337560 249300 337612
rect 249662 337900 249714 337952
rect 249754 337900 249806 337952
rect 249846 337900 249898 337952
rect 250030 337900 250082 337952
rect 250122 337900 250174 337952
rect 250214 337900 250266 337952
rect 250766 337900 250818 337952
rect 250858 337900 250910 337952
rect 251042 337900 251094 337952
rect 251410 337900 251462 337952
rect 251686 337900 251738 337952
rect 252054 337900 252106 337952
rect 252330 337900 252382 337952
rect 249478 337764 249530 337816
rect 248236 337492 248288 337544
rect 249340 337492 249392 337544
rect 248144 337424 248196 337476
rect 249616 337696 249668 337748
rect 249984 337764 250036 337816
rect 249708 337628 249760 337680
rect 249524 337560 249576 337612
rect 250582 337832 250634 337884
rect 250214 337764 250266 337816
rect 250536 337560 250588 337612
rect 250720 337560 250772 337612
rect 249892 337492 249944 337544
rect 251134 337832 251186 337884
rect 251318 337832 251370 337884
rect 251180 337696 251232 337748
rect 250996 337628 251048 337680
rect 251088 337560 251140 337612
rect 251870 337832 251922 337884
rect 251640 337764 251692 337816
rect 252238 337832 252290 337884
rect 252008 337764 252060 337816
rect 251364 337560 251416 337612
rect 251548 337560 251600 337612
rect 251732 337560 251784 337612
rect 252376 337628 252428 337680
rect 251456 337492 251508 337544
rect 252606 337832 252658 337884
rect 253434 337900 253486 337952
rect 253894 337900 253946 337952
rect 254906 337900 254958 337952
rect 255090 337900 255142 337952
rect 255182 337900 255234 337952
rect 255274 337900 255326 337952
rect 255366 337900 255418 337952
rect 253158 337832 253210 337884
rect 253250 337832 253302 337884
rect 253618 337832 253670 337884
rect 253112 337628 253164 337680
rect 253296 337628 253348 337680
rect 254262 337832 254314 337884
rect 254446 337832 254498 337884
rect 254078 337764 254130 337816
rect 253940 337696 253992 337748
rect 254216 337696 254268 337748
rect 254124 337628 254176 337680
rect 254538 337764 254590 337816
rect 254630 337764 254682 337816
rect 254722 337764 254774 337816
rect 255044 337764 255096 337816
rect 255136 337764 255188 337816
rect 252560 337560 252612 337612
rect 252836 337560 252888 337612
rect 254308 337560 254360 337612
rect 255228 337696 255280 337748
rect 254768 337628 254820 337680
rect 256194 337900 256246 337952
rect 255504 337628 255556 337680
rect 254676 337560 254728 337612
rect 255320 337560 255372 337612
rect 254492 337492 254544 337544
rect 257298 337900 257350 337952
rect 257390 337900 257442 337952
rect 257574 337900 257626 337952
rect 257942 337900 257994 337952
rect 250352 337424 250404 337476
rect 250904 337424 250956 337476
rect 256424 337492 256476 337544
rect 139400 337356 139452 337408
rect 255688 337424 255740 337476
rect 256654 337832 256706 337884
rect 256838 337832 256890 337884
rect 256792 337560 256844 337612
rect 257436 337696 257488 337748
rect 257344 337560 257396 337612
rect 257666 337832 257718 337884
rect 256976 337424 257028 337476
rect 81440 337288 81492 337340
rect 256884 337356 256936 337408
rect 257850 337764 257902 337816
rect 257804 337628 257856 337680
rect 258126 337764 258178 337816
rect 258080 337628 258132 337680
rect 257896 337560 257948 337612
rect 258402 337900 258454 337952
rect 258494 337900 258546 337952
rect 258678 337900 258730 337952
rect 258862 337900 258914 337952
rect 258954 337900 259006 337952
rect 259230 337900 259282 337952
rect 259414 337900 259466 337952
rect 259506 337900 259558 337952
rect 259598 337900 259650 337952
rect 259874 337900 259926 337952
rect 259966 337900 260018 337952
rect 260242 337900 260294 337952
rect 260426 337900 260478 337952
rect 260518 337900 260570 337952
rect 261254 337900 261306 337952
rect 261622 337900 261674 337952
rect 261714 337900 261766 337952
rect 262082 337900 262134 337952
rect 262266 337900 262318 337952
rect 262726 337900 262778 337952
rect 258448 337764 258500 337816
rect 258356 337628 258408 337680
rect 258816 337560 258868 337612
rect 259000 337560 259052 337612
rect 258264 337492 258316 337544
rect 258540 337492 258592 337544
rect 259460 337764 259512 337816
rect 259690 337832 259742 337884
rect 259552 337696 259604 337748
rect 259368 337628 259420 337680
rect 259874 337764 259926 337816
rect 259644 337492 259696 337544
rect 259828 337424 259880 337476
rect 260196 337628 260248 337680
rect 261162 337832 261214 337884
rect 260702 337764 260754 337816
rect 260564 337492 260616 337544
rect 261208 337696 261260 337748
rect 261116 337560 261168 337612
rect 262174 337832 262226 337884
rect 262036 337764 262088 337816
rect 261668 337628 261720 337680
rect 261944 337560 261996 337612
rect 261208 337492 261260 337544
rect 262450 337764 262502 337816
rect 262220 337696 262272 337748
rect 262588 337560 262640 337612
rect 262496 337492 262548 337544
rect 260472 337424 260524 337476
rect 260656 337424 260708 337476
rect 259920 337356 259972 337408
rect 262910 337900 262962 337952
rect 263002 337900 263054 337952
rect 263094 337900 263146 337952
rect 263554 337900 263606 337952
rect 263646 337900 263698 337952
rect 264014 337900 264066 337952
rect 265486 337900 265538 337952
rect 262956 337764 263008 337816
rect 263278 337764 263330 337816
rect 263140 337628 263192 337680
rect 263232 337424 263284 337476
rect 263508 337424 263560 337476
rect 263830 337832 263882 337884
rect 263876 337696 263928 337748
rect 264658 337832 264710 337884
rect 264750 337832 264802 337884
rect 265026 337832 265078 337884
rect 265302 337832 265354 337884
rect 264198 337764 264250 337816
rect 264382 337764 264434 337816
rect 264060 337628 264112 337680
rect 263692 337424 263744 337476
rect 264428 337628 264480 337680
rect 264244 337356 264296 337408
rect 26240 337220 26292 337272
rect 242992 337220 243044 337272
rect 248972 337288 249024 337340
rect 253940 337288 253992 337340
rect 264152 337288 264204 337340
rect 264612 337492 264664 337544
rect 265072 337696 265124 337748
rect 265348 337696 265400 337748
rect 265164 337492 265216 337544
rect 265670 337832 265722 337884
rect 265716 337696 265768 337748
rect 265624 337628 265676 337680
rect 265716 337560 265768 337612
rect 264980 337424 265032 337476
rect 266958 337900 267010 337952
rect 267050 337900 267102 337952
rect 267142 337900 267194 337952
rect 267510 337900 267562 337952
rect 268062 337900 268114 337952
rect 269074 337900 269126 337952
rect 269350 337900 269402 337952
rect 269718 337900 269770 337952
rect 269810 337900 269862 337952
rect 265946 337832 265998 337884
rect 266498 337832 266550 337884
rect 266590 337832 266642 337884
rect 266084 337560 266136 337612
rect 265900 337424 265952 337476
rect 265808 337356 265860 337408
rect 267004 337764 267056 337816
rect 267234 337832 267286 337884
rect 267326 337832 267378 337884
rect 266636 337696 266688 337748
rect 267096 337696 267148 337748
rect 267188 337628 267240 337680
rect 267464 337628 267516 337680
rect 267372 337560 267424 337612
rect 268338 337832 268390 337884
rect 268798 337832 268850 337884
rect 266636 337492 266688 337544
rect 267740 337492 267792 337544
rect 268476 337492 268528 337544
rect 268108 337424 268160 337476
rect 268936 337628 268988 337680
rect 269166 337832 269218 337884
rect 269304 337628 269356 337680
rect 270086 337832 270138 337884
rect 269534 337764 269586 337816
rect 269764 337764 269816 337816
rect 269488 337628 269540 337680
rect 269580 337628 269632 337680
rect 270040 337560 270092 337612
rect 270270 337900 270322 337952
rect 270362 337900 270414 337952
rect 270730 337900 270782 337952
rect 271098 337900 271150 337952
rect 271190 337900 271242 337952
rect 270408 337764 270460 337816
rect 270914 337832 270966 337884
rect 270776 337560 270828 337612
rect 269212 337492 269264 337544
rect 270592 337492 270644 337544
rect 271558 337832 271610 337884
rect 271834 337832 271886 337884
rect 271236 337628 271288 337680
rect 271696 337628 271748 337680
rect 272202 337900 272254 337952
rect 272570 337900 272622 337952
rect 272938 337900 272990 337952
rect 273122 337900 273174 337952
rect 273766 337900 273818 337952
rect 274134 337900 274186 337952
rect 274226 337900 274278 337952
rect 274318 337900 274370 337952
rect 274502 337900 274554 337952
rect 272432 337628 272484 337680
rect 272524 337628 272576 337680
rect 272984 337628 273036 337680
rect 272340 337560 272392 337612
rect 271972 337492 272024 337544
rect 273306 337832 273358 337884
rect 273490 337832 273542 337884
rect 273950 337832 274002 337884
rect 274042 337832 274094 337884
rect 273720 337764 273772 337816
rect 273628 337628 273680 337680
rect 274134 337764 274186 337816
rect 274364 337764 274416 337816
rect 274456 337764 274508 337816
rect 274548 337696 274600 337748
rect 274778 337764 274830 337816
rect 274088 337560 274140 337612
rect 274272 337560 274324 337612
rect 273996 337492 274048 337544
rect 274180 337492 274232 337544
rect 274962 337900 275014 337952
rect 275054 337832 275106 337884
rect 275146 337832 275198 337884
rect 275008 337628 275060 337680
rect 275514 337900 275566 337952
rect 275606 337832 275658 337884
rect 275560 337696 275612 337748
rect 275882 337900 275934 337952
rect 276158 337900 276210 337952
rect 276250 337900 276302 337952
rect 276342 337900 276394 337952
rect 276526 337900 276578 337952
rect 276618 337900 276670 337952
rect 276802 337900 276854 337952
rect 276894 337900 276946 337952
rect 276986 337900 277038 337952
rect 275468 337628 275520 337680
rect 275744 337628 275796 337680
rect 274824 337424 274876 337476
rect 274732 337356 274784 337408
rect 251640 337220 251692 337272
rect 275376 337560 275428 337612
rect 275974 337832 276026 337884
rect 276204 337764 276256 337816
rect 276296 337628 276348 337680
rect 276020 337560 276072 337612
rect 276664 337628 276716 337680
rect 276572 337492 276624 337544
rect 276388 337424 276440 337476
rect 276848 337764 276900 337816
rect 276940 337696 276992 337748
rect 277262 337900 277314 337952
rect 277630 337900 277682 337952
rect 277814 337900 277866 337952
rect 277906 337900 277958 337952
rect 277998 337900 278050 337952
rect 278090 337900 278142 337952
rect 278182 337900 278234 337952
rect 277032 337628 277084 337680
rect 277124 337492 277176 337544
rect 277676 337628 277728 337680
rect 278044 337764 278096 337816
rect 277952 337560 278004 337612
rect 277860 337492 277912 337544
rect 278366 337764 278418 337816
rect 278734 337900 278786 337952
rect 278918 337900 278970 337952
rect 279010 337900 279062 337952
rect 279102 337900 279154 337952
rect 279194 337900 279246 337952
rect 279286 337900 279338 337952
rect 278780 337764 278832 337816
rect 278964 337696 279016 337748
rect 278320 337628 278372 337680
rect 278596 337628 278648 337680
rect 278688 337628 278740 337680
rect 278872 337560 278924 337612
rect 279470 337900 279522 337952
rect 279562 337900 279614 337952
rect 279654 337900 279706 337952
rect 279838 337900 279890 337952
rect 280022 337900 280074 337952
rect 279240 337560 279292 337612
rect 279332 337560 279384 337612
rect 279148 337492 279200 337544
rect 278136 337424 278188 337476
rect 279516 337696 279568 337748
rect 279608 337696 279660 337748
rect 279792 337492 279844 337544
rect 279976 337764 280028 337816
rect 430580 338240 430632 338292
rect 448520 338172 448572 338224
rect 280206 337900 280258 337952
rect 280482 337832 280534 337884
rect 280574 337832 280626 337884
rect 280528 337628 280580 337680
rect 280344 337560 280396 337612
rect 280436 337560 280488 337612
rect 281034 337900 281086 337952
rect 281402 337900 281454 337952
rect 280942 337832 280994 337884
rect 281126 337832 281178 337884
rect 281310 337832 281362 337884
rect 281218 337764 281270 337816
rect 281080 337696 281132 337748
rect 280988 337560 281040 337612
rect 281172 337560 281224 337612
rect 281264 337492 281316 337544
rect 279884 337424 279936 337476
rect 280804 337424 280856 337476
rect 465080 338104 465132 338156
rect 290924 338036 290976 338088
rect 281770 337900 281822 337952
rect 282138 337900 282190 337952
rect 282230 337900 282282 337952
rect 282966 337900 283018 337952
rect 283978 337900 284030 337952
rect 284346 337900 284398 337952
rect 284530 337900 284582 337952
rect 281586 337832 281638 337884
rect 281954 337832 282006 337884
rect 281540 337628 281592 337680
rect 281632 337560 281684 337612
rect 282092 337696 282144 337748
rect 282598 337832 282650 337884
rect 282874 337832 282926 337884
rect 282276 337628 282328 337680
rect 282644 337560 282696 337612
rect 280068 337356 280120 337408
rect 281448 337356 281500 337408
rect 275192 337288 275244 337340
rect 282460 337288 282512 337340
rect 275100 337220 275152 337272
rect 280252 337220 280304 337272
rect 281448 337220 281500 337272
rect 281908 337220 281960 337272
rect 283334 337832 283386 337884
rect 283610 337832 283662 337884
rect 283150 337764 283202 337816
rect 283104 337628 283156 337680
rect 283932 337764 283984 337816
rect 284070 337764 284122 337816
rect 284254 337764 284306 337816
rect 284024 337628 284076 337680
rect 284622 337832 284674 337884
rect 284714 337832 284766 337884
rect 284484 337696 284536 337748
rect 284576 337628 284628 337680
rect 284392 337560 284444 337612
rect 284668 337560 284720 337612
rect 283288 337492 283340 337544
rect 283472 337492 283524 337544
rect 284208 337492 284260 337544
rect 285266 337900 285318 337952
rect 286462 337900 286514 337952
rect 286554 337900 286606 337952
rect 286646 337900 286698 337952
rect 287014 337900 287066 337952
rect 287198 337900 287250 337952
rect 287382 337900 287434 337952
rect 287566 337900 287618 337952
rect 287658 337900 287710 337952
rect 287934 337900 287986 337952
rect 288026 337900 288078 337952
rect 288210 337900 288262 337952
rect 288578 337900 288630 337952
rect 289222 337900 289274 337952
rect 289682 337900 289734 337952
rect 285174 337832 285226 337884
rect 285358 337832 285410 337884
rect 285450 337832 285502 337884
rect 285542 337832 285594 337884
rect 286094 337832 286146 337884
rect 285312 337628 285364 337680
rect 285404 337628 285456 337680
rect 285128 337492 285180 337544
rect 285036 337424 285088 337476
rect 285220 337424 285272 337476
rect 286508 337764 286560 337816
rect 286600 337764 286652 337816
rect 286830 337764 286882 337816
rect 287244 337764 287296 337816
rect 286692 337628 286744 337680
rect 286876 337628 286928 337680
rect 286232 337560 286284 337612
rect 287520 337764 287572 337816
rect 287842 337764 287894 337816
rect 287612 337628 287664 337680
rect 287796 337628 287848 337680
rect 287704 337560 287756 337612
rect 287152 337492 287204 337544
rect 287612 337492 287664 337544
rect 286968 337424 287020 337476
rect 288302 337832 288354 337884
rect 288210 337764 288262 337816
rect 288670 337832 288722 337884
rect 288854 337764 288906 337816
rect 288624 337696 288676 337748
rect 288256 337628 288308 337680
rect 288072 337560 288124 337612
rect 288946 337696 288998 337748
rect 288808 337492 288860 337544
rect 288440 337424 288492 337476
rect 289314 337764 289366 337816
rect 289406 337764 289458 337816
rect 290832 337968 290884 338020
rect 290050 337900 290102 337952
rect 290234 337900 290286 337952
rect 290326 337900 290378 337952
rect 290510 337900 290562 337952
rect 289866 337832 289918 337884
rect 289958 337832 290010 337884
rect 289176 337628 289228 337680
rect 289636 337696 289688 337748
rect 290096 337696 290148 337748
rect 289728 337628 289780 337680
rect 289912 337628 289964 337680
rect 289084 337560 289136 337612
rect 289360 337560 289412 337612
rect 289820 337560 289872 337612
rect 290372 337628 290424 337680
rect 290464 337628 290516 337680
rect 283748 337356 283800 337408
rect 287612 337356 287664 337408
rect 346584 337356 346636 337408
rect 283564 337288 283616 337340
rect 288072 337288 288124 337340
rect 346676 337288 346728 337340
rect 283748 337220 283800 337272
rect 285588 337220 285640 337272
rect 345664 337220 345716 337272
rect 227720 337152 227772 337204
rect 263140 337152 263192 337204
rect 271880 337152 271932 337204
rect 218060 337084 218112 337136
rect 262220 337084 262272 337136
rect 346492 337152 346544 337204
rect 275744 337084 275796 337136
rect 343916 337084 343968 337136
rect 165620 337016 165672 337068
rect 248972 337016 249024 337068
rect 250168 337016 250220 337068
rect 250628 337016 250680 337068
rect 161480 336948 161532 337000
rect 257896 336948 257948 337000
rect 270040 336948 270092 337000
rect 346400 337016 346452 337068
rect 276112 336948 276164 337000
rect 394700 336948 394752 337000
rect 241428 336880 241480 336932
rect 249800 336880 249852 336932
rect 240048 336812 240100 336864
rect 267280 336880 267332 336932
rect 272432 336880 272484 336932
rect 273628 336812 273680 336864
rect 234620 336744 234672 336796
rect 263692 336744 263744 336796
rect 242348 336676 242400 336728
rect 246764 336676 246816 336728
rect 256424 336676 256476 336728
rect 268200 336676 268252 336728
rect 244188 336608 244240 336660
rect 248420 336608 248472 336660
rect 260932 336608 260984 336660
rect 277216 336880 277268 336932
rect 408500 336880 408552 336932
rect 280344 336812 280396 336864
rect 451280 336812 451332 336864
rect 280252 336744 280304 336796
rect 281172 336744 281224 336796
rect 281724 336744 281776 336796
rect 282552 336744 282604 336796
rect 292856 336744 292908 336796
rect 557540 336744 557592 336796
rect 285588 336676 285640 336728
rect 287244 336676 287296 336728
rect 291200 336676 291252 336728
rect 277308 336608 277360 336660
rect 264980 336540 265032 336592
rect 274732 336540 274784 336592
rect 287612 336608 287664 336660
rect 279792 336540 279844 336592
rect 285312 336540 285364 336592
rect 287244 336540 287296 336592
rect 293408 336540 293460 336592
rect 224960 336472 225012 336524
rect 262312 336472 262364 336524
rect 278688 336472 278740 336524
rect 287888 336472 287940 336524
rect 196624 336404 196676 336456
rect 247776 336404 247828 336456
rect 277400 336404 277452 336456
rect 293224 336404 293276 336456
rect 200764 336336 200816 336388
rect 248604 336336 248656 336388
rect 249800 336336 249852 336388
rect 188344 336268 188396 336320
rect 247500 336268 247552 336320
rect 255504 336268 255556 336320
rect 256608 336268 256660 336320
rect 258448 336268 258500 336320
rect 259184 336268 259236 336320
rect 259736 336268 259788 336320
rect 260288 336268 260340 336320
rect 182180 336200 182232 336252
rect 248972 336200 249024 336252
rect 253572 336200 253624 336252
rect 262680 336200 262732 336252
rect 276020 336336 276072 336388
rect 291936 336336 291988 336388
rect 280712 336268 280764 336320
rect 346768 336268 346820 336320
rect 266268 336200 266320 336252
rect 270408 336200 270460 336252
rect 279884 336200 279936 336252
rect 281540 336200 281592 336252
rect 467840 336200 467892 336252
rect 160100 336132 160152 336184
rect 257804 336132 257856 336184
rect 257896 336132 257948 336184
rect 264244 336132 264296 336184
rect 277584 336132 277636 336184
rect 278964 336132 279016 336184
rect 281356 336132 281408 336184
rect 283196 336132 283248 336184
rect 283748 336132 283800 336184
rect 483020 336132 483072 336184
rect 128360 336064 128412 336116
rect 255320 336064 255372 336116
rect 125600 335996 125652 336048
rect 255044 335996 255096 336048
rect 242440 335928 242492 335980
rect 253296 335928 253348 335980
rect 255320 335928 255372 335980
rect 267740 336064 267792 336116
rect 281540 336064 281592 336116
rect 282276 336064 282328 336116
rect 284392 336064 284444 336116
rect 500960 336064 501012 336116
rect 256424 335996 256476 336048
rect 273260 335996 273312 336048
rect 287060 335996 287112 336048
rect 536840 335996 536892 336048
rect 259184 335928 259236 335980
rect 268476 335928 268528 335980
rect 269948 335928 270000 335980
rect 270224 335928 270276 335980
rect 278136 335928 278188 335980
rect 292120 335928 292172 335980
rect 243728 335860 243780 335912
rect 251916 335860 251968 335912
rect 260012 335860 260064 335912
rect 260288 335860 260340 335912
rect 262680 335860 262732 335912
rect 262956 335860 263008 335912
rect 277400 335860 277452 335912
rect 277768 335860 277820 335912
rect 278596 335860 278648 335912
rect 287244 335860 287296 335912
rect 287888 335860 287940 335912
rect 293316 335860 293368 335912
rect 242164 335792 242216 335844
rect 248420 335792 248472 335844
rect 248972 335792 249024 335844
rect 259460 335792 259512 335844
rect 279332 335792 279384 335844
rect 293500 335792 293552 335844
rect 243912 335724 243964 335776
rect 252468 335724 252520 335776
rect 255780 335724 255832 335776
rect 255964 335724 256016 335776
rect 261300 335724 261352 335776
rect 261576 335724 261628 335776
rect 283196 335724 283248 335776
rect 294604 335724 294656 335776
rect 248972 335656 249024 335708
rect 261760 335656 261812 335708
rect 273168 335656 273220 335708
rect 288072 335656 288124 335708
rect 251916 335588 251968 335640
rect 255872 335588 255924 335640
rect 277308 335588 277360 335640
rect 281356 335588 281408 335640
rect 252468 335520 252520 335572
rect 261576 335520 261628 335572
rect 265348 335520 265400 335572
rect 276204 335520 276256 335572
rect 292028 335588 292080 335640
rect 258172 335452 258224 335504
rect 274916 335452 274968 335504
rect 281816 335452 281868 335504
rect 252192 335384 252244 335436
rect 258356 335384 258408 335436
rect 274824 335384 274876 335436
rect 275008 335384 275060 335436
rect 276112 335384 276164 335436
rect 276664 335384 276716 335436
rect 254492 335316 254544 335368
rect 260840 335316 260892 335368
rect 274732 335316 274784 335368
rect 275376 335316 275428 335368
rect 275836 335316 275888 335368
rect 283748 335316 283800 335368
rect 285680 335316 285732 335368
rect 286416 335316 286468 335368
rect 288348 335316 288400 335368
rect 291844 335316 291896 335368
rect 255688 335248 255740 335300
rect 256332 335248 256384 335300
rect 272340 335248 272392 335300
rect 346860 335248 346912 335300
rect 242900 335180 242952 335232
rect 257896 335180 257948 335232
rect 274272 335180 274324 335232
rect 349160 335180 349212 335232
rect 242256 335112 242308 335164
rect 259920 335112 259972 335164
rect 272708 335112 272760 335164
rect 351920 335112 351972 335164
rect 233240 335044 233292 335096
rect 263416 335044 263468 335096
rect 283472 335044 283524 335096
rect 491300 335044 491352 335096
rect 229100 334976 229152 335028
rect 263048 334976 263100 335028
rect 285588 334976 285640 335028
rect 509240 334976 509292 335028
rect 211160 334908 211212 334960
rect 248972 334908 249024 334960
rect 249248 334908 249300 334960
rect 249432 334908 249484 334960
rect 173900 334840 173952 334892
rect 258816 334908 258868 334960
rect 274548 334908 274600 334960
rect 279884 334908 279936 334960
rect 286232 334908 286284 334960
rect 523040 334908 523092 334960
rect 151820 334772 151872 334824
rect 257160 334840 257212 334892
rect 286692 334840 286744 334892
rect 531320 334840 531372 334892
rect 136640 334704 136692 334756
rect 256056 334772 256108 334824
rect 290924 334772 290976 334824
rect 538220 334772 538272 334824
rect 133880 334636 133932 334688
rect 255964 334704 256016 334756
rect 291016 334704 291068 334756
rect 545120 334704 545172 334756
rect 288624 334636 288676 334688
rect 556160 334636 556212 334688
rect 249248 334568 249300 334620
rect 251364 334568 251416 334620
rect 253204 334568 253256 334620
rect 253480 334568 253532 334620
rect 253940 334568 253992 334620
rect 255136 334568 255188 334620
rect 264244 334568 264296 334620
rect 264612 334568 264664 334620
rect 265440 334568 265492 334620
rect 265808 334568 265860 334620
rect 266728 334568 266780 334620
rect 267188 334568 267240 334620
rect 283196 334568 283248 334620
rect 283380 334568 283432 334620
rect 284392 334568 284444 334620
rect 284852 334568 284904 334620
rect 289636 334568 289688 334620
rect 565820 334568 565872 334620
rect 52460 334500 52512 334552
rect 247040 334500 247092 334552
rect 248880 334500 248932 334552
rect 249156 334500 249208 334552
rect 273812 334432 273864 334484
rect 276756 334432 276808 334484
rect 249156 334364 249208 334416
rect 259000 334364 259052 334416
rect 288532 334364 288584 334416
rect 289360 334364 289412 334416
rect 265716 334228 265768 334280
rect 266268 334228 266320 334280
rect 285772 334024 285824 334076
rect 286600 334024 286652 334076
rect 149060 333820 149112 333872
rect 256700 333820 256752 333872
rect 241520 333752 241572 333804
rect 216680 333684 216732 333736
rect 261208 333752 261260 333804
rect 263968 333752 264020 333804
rect 155960 333616 156012 333668
rect 257528 333616 257580 333668
rect 255320 333548 255372 333600
rect 256424 333548 256476 333600
rect 257436 333548 257488 333600
rect 301136 333548 301188 333600
rect 135260 333480 135312 333532
rect 255596 333480 255648 333532
rect 276480 333480 276532 333532
rect 398840 333480 398892 333532
rect 118700 333412 118752 333464
rect 254584 333412 254636 333464
rect 265624 333412 265676 333464
rect 276940 333412 276992 333464
rect 407120 333412 407172 333464
rect 91100 333344 91152 333396
rect 252284 333344 252336 333396
rect 256240 333344 256292 333396
rect 273812 333344 273864 333396
rect 274180 333344 274232 333396
rect 278964 333344 279016 333396
rect 414020 333344 414072 333396
rect 84200 333276 84252 333328
rect 251548 333276 251600 333328
rect 279148 333276 279200 333328
rect 420920 333276 420972 333328
rect 41420 333208 41472 333260
rect 245384 333208 245436 333260
rect 247132 333208 247184 333260
rect 248052 333208 248104 333260
rect 250076 333208 250128 333260
rect 250260 333208 250312 333260
rect 250352 333208 250404 333260
rect 250720 333208 250772 333260
rect 271972 333208 272024 333260
rect 272248 333208 272300 333260
rect 272524 333208 272576 333260
rect 274180 333208 274232 333260
rect 277584 333208 277636 333260
rect 278320 333208 278372 333260
rect 280068 333208 280120 333260
rect 438860 333208 438912 333260
rect 247776 333140 247828 333192
rect 248788 333140 248840 333192
rect 249984 333140 250036 333192
rect 250812 333140 250864 333192
rect 274364 333140 274416 333192
rect 276572 333140 276624 333192
rect 248696 333072 248748 333124
rect 249432 333072 249484 333124
rect 250260 333072 250312 333124
rect 250996 333072 251048 333124
rect 247408 333004 247460 333056
rect 247960 333004 248012 333056
rect 248788 333004 248840 333056
rect 249616 333004 249668 333056
rect 272432 333004 272484 333056
rect 272616 333004 272668 333056
rect 246764 332936 246816 332988
rect 265808 332936 265860 332988
rect 273536 332868 273588 332920
rect 274088 332868 274140 332920
rect 243636 332324 243688 332376
rect 260748 332324 260800 332376
rect 226340 332256 226392 332308
rect 262680 332256 262732 332308
rect 233884 332188 233936 332240
rect 258540 332188 258592 332240
rect 259920 332188 259972 332240
rect 300952 332188 301004 332240
rect 257804 332120 257856 332172
rect 301044 332120 301096 332172
rect 168380 332052 168432 332104
rect 246856 332052 246908 332104
rect 272984 332052 273036 332104
rect 354680 332052 354732 332104
rect 122840 331984 122892 332036
rect 255412 331984 255464 332036
rect 281816 331984 281868 332036
rect 379520 331984 379572 332036
rect 74540 331916 74592 331968
rect 251180 331916 251232 331968
rect 289084 331916 289136 331968
rect 556252 331916 556304 331968
rect 34520 331848 34572 331900
rect 247592 331848 247644 331900
rect 289176 331848 289228 331900
rect 564440 331848 564492 331900
rect 248972 331644 249024 331696
rect 249708 331644 249760 331696
rect 260748 331236 260800 331288
rect 265992 331236 266044 331288
rect 257252 331168 257304 331220
rect 257528 331168 257580 331220
rect 251640 330964 251692 331016
rect 251916 330964 251968 331016
rect 272156 330964 272208 331016
rect 272800 330964 272852 331016
rect 251180 330896 251232 330948
rect 252468 330896 252520 330948
rect 234712 330828 234764 330880
rect 263416 330828 263468 330880
rect 207020 330760 207072 330812
rect 261300 330760 261352 330812
rect 266452 330760 266504 330812
rect 269120 330760 269172 330812
rect 270224 330760 270276 330812
rect 193220 330692 193272 330744
rect 259552 330692 259604 330744
rect 184940 330624 184992 330676
rect 251180 330624 251232 330676
rect 251364 330624 251416 330676
rect 252008 330624 252060 330676
rect 252836 330624 252888 330676
rect 253112 330624 253164 330676
rect 255964 330624 256016 330676
rect 264888 330692 264940 330744
rect 263784 330624 263836 330676
rect 264336 330624 264388 330676
rect 189080 330556 189132 330608
rect 260288 330556 260340 330608
rect 263968 330556 264020 330608
rect 264796 330556 264848 330608
rect 269304 330692 269356 330744
rect 270040 330692 270092 330744
rect 266912 330624 266964 330676
rect 266544 330556 266596 330608
rect 60740 330488 60792 330540
rect 245752 330488 245804 330540
rect 245844 330488 245896 330540
rect 246580 330488 246632 330540
rect 247868 330488 247920 330540
rect 248328 330488 248380 330540
rect 251548 330488 251600 330540
rect 252100 330488 252152 330540
rect 252560 330488 252612 330540
rect 252836 330488 252888 330540
rect 253296 330488 253348 330540
rect 253756 330488 253808 330540
rect 264060 330488 264112 330540
rect 264336 330488 264388 330540
rect 265256 330488 265308 330540
rect 265532 330488 265584 330540
rect 269120 330624 269172 330676
rect 269580 330624 269632 330676
rect 268292 330488 268344 330540
rect 268476 330488 268528 330540
rect 269580 330488 269632 330540
rect 269856 330488 269908 330540
rect 271144 330624 271196 330676
rect 281356 330624 281408 330676
rect 361580 330624 361632 330676
rect 275652 330556 275704 330608
rect 358820 330556 358872 330608
rect 290832 330488 290884 330540
rect 572720 330488 572772 330540
rect 246120 330420 246172 330472
rect 246672 330420 246724 330472
rect 251456 330420 251508 330472
rect 252376 330420 252428 330472
rect 253020 330420 253072 330472
rect 253848 330420 253900 330472
rect 263876 330420 263928 330472
rect 264428 330420 264480 330472
rect 267004 330420 267056 330472
rect 268016 330420 268068 330472
rect 268200 330420 268252 330472
rect 269212 330420 269264 330472
rect 269396 330420 269448 330472
rect 269488 330420 269540 330472
rect 269948 330420 270000 330472
rect 271052 330420 271104 330472
rect 245752 330352 245804 330404
rect 246948 330352 247000 330404
rect 252652 330352 252704 330404
rect 253664 330352 253716 330404
rect 264060 330352 264112 330404
rect 264520 330352 264572 330404
rect 265532 330352 265584 330404
rect 266084 330352 266136 330404
rect 266728 330352 266780 330404
rect 267372 330352 267424 330404
rect 268292 330352 268344 330404
rect 268568 330352 268620 330404
rect 270868 330352 270920 330404
rect 271328 330352 271380 330404
rect 251640 330284 251692 330336
rect 251824 330284 251876 330336
rect 254952 330284 255004 330336
rect 264612 330284 264664 330336
rect 268200 330284 268252 330336
rect 268752 330284 268804 330336
rect 269396 330284 269448 330336
rect 270132 330284 270184 330336
rect 270684 330284 270736 330336
rect 271604 330284 271656 330336
rect 267740 330216 267792 330268
rect 268568 330216 268620 330268
rect 265348 329672 265400 329724
rect 266176 329672 266228 329724
rect 220820 329332 220872 329384
rect 253480 329332 253532 329384
rect 153200 329264 153252 329316
rect 256976 329264 257028 329316
rect 126980 329196 127032 329248
rect 253940 329196 253992 329248
rect 52552 329128 52604 329180
rect 248144 329128 248196 329180
rect 283656 329128 283708 329180
rect 489920 329128 489972 329180
rect 37280 329060 37332 329112
rect 248236 329060 248288 329112
rect 287612 329060 287664 329112
rect 539600 329060 539652 329112
rect 283012 328380 283064 328432
rect 283472 328380 283524 328432
rect 274640 328108 274692 328160
rect 275652 328108 275704 328160
rect 180800 327836 180852 327888
rect 259368 327836 259420 327888
rect 276940 327836 276992 327888
rect 398932 327836 398984 327888
rect 171140 327768 171192 327820
rect 252192 327768 252244 327820
rect 278228 327768 278280 327820
rect 423680 327768 423732 327820
rect 46940 327700 46992 327752
rect 249064 327700 249116 327752
rect 290188 327700 290240 327752
rect 575480 327700 575532 327752
rect 276296 327360 276348 327412
rect 276940 327360 276992 327412
rect 285128 326748 285180 326800
rect 294512 326748 294564 326800
rect 257160 326680 257212 326732
rect 257988 326680 258040 326732
rect 274732 326680 274784 326732
rect 284300 326680 284352 326732
rect 285312 326680 285364 326732
rect 257620 326544 257672 326596
rect 257988 326544 258040 326596
rect 261392 326544 261444 326596
rect 261760 326544 261812 326596
rect 209780 326340 209832 326392
rect 261944 326476 261996 326528
rect 279884 326612 279936 326664
rect 288624 326612 288676 326664
rect 288808 326612 288860 326664
rect 365720 326612 365772 326664
rect 275284 326544 275336 326596
rect 286048 326544 286100 326596
rect 254308 326408 254360 326460
rect 254768 326408 254820 326460
rect 256148 326408 256200 326460
rect 256516 326408 256568 326460
rect 262496 326408 262548 326460
rect 263232 326408 263284 326460
rect 274732 326408 274784 326460
rect 254492 326340 254544 326392
rect 255228 326340 255280 326392
rect 256976 326340 257028 326392
rect 257712 326340 257764 326392
rect 258264 326340 258316 326392
rect 259276 326340 259328 326392
rect 260012 326340 260064 326392
rect 260656 326340 260708 326392
rect 261300 326340 261352 326392
rect 261852 326340 261904 326392
rect 262680 326340 262732 326392
rect 263324 326340 263376 326392
rect 275192 326340 275244 326392
rect 286416 326476 286468 326528
rect 294512 326544 294564 326596
rect 512000 326544 512052 326596
rect 277584 326408 277636 326460
rect 277676 326408 277728 326460
rect 277860 326408 277912 326460
rect 282000 326408 282052 326460
rect 282276 326408 282328 326460
rect 284484 326408 284536 326460
rect 284852 326408 284904 326460
rect 289912 326408 289964 326460
rect 523132 326476 523184 326528
rect 528560 326408 528612 326460
rect 276020 326340 276072 326392
rect 276848 326340 276900 326392
rect 254216 326272 254268 326324
rect 254860 326272 254912 326324
rect 261392 326272 261444 326324
rect 262036 326272 262088 326324
rect 278964 326340 279016 326392
rect 279608 326340 279660 326392
rect 280528 326340 280580 326392
rect 281264 326340 281316 326392
rect 287244 326340 287296 326392
rect 287428 326340 287480 326392
rect 288808 326340 288860 326392
rect 289452 326340 289504 326392
rect 572812 326340 572864 326392
rect 280620 326272 280672 326324
rect 280804 326272 280856 326324
rect 256332 326204 256384 326256
rect 260196 326204 260248 326256
rect 260380 326204 260432 326256
rect 275284 326204 275336 326256
rect 275560 326204 275612 326256
rect 276296 326204 276348 326256
rect 276664 326204 276716 326256
rect 277768 326204 277820 326256
rect 284576 326204 284628 326256
rect 284760 326204 284812 326256
rect 285956 326204 286008 326256
rect 286140 326204 286192 326256
rect 287428 326204 287480 326256
rect 287796 326204 287848 326256
rect 289820 326204 289872 326256
rect 290740 326204 290792 326256
rect 254676 325932 254728 325984
rect 254952 325932 255004 325984
rect 258448 326136 258500 326188
rect 259000 326136 259052 326188
rect 274916 326136 274968 326188
rect 275468 326136 275520 326188
rect 277492 326136 277544 326188
rect 278136 326136 278188 326188
rect 275008 326068 275060 326120
rect 275836 326068 275888 326120
rect 284760 326068 284812 326120
rect 285036 326068 285088 326120
rect 285680 326068 285732 326120
rect 285956 326068 286008 326120
rect 256424 325932 256476 325984
rect 273352 325864 273404 325916
rect 273904 325864 273956 325916
rect 279056 325796 279108 325848
rect 279332 325796 279384 325848
rect 279516 325728 279568 325780
rect 278780 325524 278832 325576
rect 279424 325524 279476 325576
rect 278780 325388 278832 325440
rect 275652 324980 275704 325032
rect 376760 324980 376812 325032
rect 280896 324912 280948 324964
rect 456800 324912 456852 324964
rect 259736 324164 259788 324216
rect 260564 324164 260616 324216
rect 20 323552 72 323604
rect 244832 323552 244884 323604
rect 276940 323552 276992 323604
rect 396080 323552 396132 323604
rect 258540 323008 258592 323060
rect 258724 323008 258776 323060
rect 261024 323008 261076 323060
rect 262128 323008 262180 323060
rect 281816 322600 281868 322652
rect 282552 322600 282604 322652
rect 191840 320832 191892 320884
rect 260196 320832 260248 320884
rect 523684 320832 523736 320884
rect 580264 320832 580316 320884
rect 247132 320764 247184 320816
rect 247316 320764 247368 320816
rect 3148 320084 3200 320136
rect 235448 320152 235500 320204
rect 245108 320152 245160 320204
rect 578148 313216 578200 313268
rect 580080 313216 580132 313268
rect 3332 306280 3384 306332
rect 233792 306280 233844 306332
rect 301872 302880 301924 302932
rect 345112 302880 345164 302932
rect 3240 293904 3292 293956
rect 235356 293904 235408 293956
rect 578056 273164 578108 273216
rect 580080 273164 580132 273216
rect 3332 266976 3384 267028
rect 232504 266976 232556 267028
rect 300492 262828 300544 262880
rect 345204 262828 345256 262880
rect 290740 260108 290792 260160
rect 443000 260108 443052 260160
rect 577964 259360 578016 259412
rect 580080 259360 580132 259412
rect 3332 255212 3384 255264
rect 91744 255212 91796 255264
rect 3332 241408 3384 241460
rect 90456 241408 90508 241460
rect 577780 219172 577832 219224
rect 579712 219172 579764 219224
rect 3332 214548 3384 214600
rect 237472 214548 237524 214600
rect 287612 193808 287664 193860
rect 547880 193808 547932 193860
rect 154580 191088 154632 191140
rect 257068 191088 257120 191140
rect 294604 184220 294656 184272
rect 449900 184220 449952 184272
rect 282184 184152 282236 184204
rect 471980 184152 472032 184204
rect 277952 180140 278004 180192
rect 418160 180140 418212 180192
rect 290188 180072 290240 180124
rect 581000 180072 581052 180124
rect 577872 179324 577924 179376
rect 579712 179324 579764 179376
rect 160192 179120 160244 179172
rect 256976 179120 257028 179172
rect 115940 179052 115992 179104
rect 254400 179052 254452 179104
rect 273812 179052 273864 179104
rect 368480 179052 368532 179104
rect 109040 178984 109092 179036
rect 253296 178984 253348 179036
rect 283564 178984 283616 179036
rect 386420 178984 386472 179036
rect 104900 178916 104952 178968
rect 253204 178916 253256 178968
rect 277860 178916 277912 178968
rect 415400 178916 415452 178968
rect 98000 178848 98052 178900
rect 253112 178848 253164 178900
rect 288900 178848 288952 178900
rect 560300 178848 560352 178900
rect 67640 178780 67692 178832
rect 250536 178780 250588 178832
rect 288808 178780 288860 178832
rect 567200 178780 567252 178832
rect 49700 178712 49752 178764
rect 248880 178712 248932 178764
rect 290004 178712 290056 178764
rect 574100 178712 574152 178764
rect 2780 178644 2832 178696
rect 244464 178644 244516 178696
rect 290096 178644 290148 178696
rect 578240 178644 578292 178696
rect 176660 177828 176712 177880
rect 258448 177828 258500 177880
rect 162860 177760 162912 177812
rect 257160 177760 257212 177812
rect 280712 177760 280764 177812
rect 452660 177760 452712 177812
rect 158720 177692 158772 177744
rect 256884 177692 256936 177744
rect 280804 177692 280856 177744
rect 459560 177692 459612 177744
rect 151912 177624 151964 177676
rect 257436 177624 257488 177676
rect 284852 177624 284904 177676
rect 503720 177624 503772 177676
rect 144920 177556 144972 177608
rect 255688 177556 255740 177608
rect 284944 177556 284996 177608
rect 510620 177556 510672 177608
rect 66260 177488 66312 177540
rect 250444 177488 250496 177540
rect 286140 177488 286192 177540
rect 521660 177488 521712 177540
rect 55220 177420 55272 177472
rect 248788 177420 248840 177472
rect 286048 177420 286100 177472
rect 524420 177420 524472 177472
rect 48320 177352 48372 177404
rect 248696 177352 248748 177404
rect 287520 177352 287572 177404
rect 542360 177352 542412 177404
rect 17960 177284 18012 177336
rect 246120 177284 246172 177336
rect 287428 177284 287480 177336
rect 546500 177284 546552 177336
rect 275376 176400 275428 176452
rect 382280 176400 382332 176452
rect 275192 176332 275244 176384
rect 385040 176332 385092 176384
rect 275284 176264 275336 176316
rect 389180 176264 389232 176316
rect 276296 176196 276348 176248
rect 402980 176196 403032 176248
rect 277676 176128 277728 176180
rect 416780 176128 416832 176180
rect 293500 176060 293552 176112
rect 436100 176060 436152 176112
rect 277768 175992 277820 176044
rect 423772 175992 423824 176044
rect 279424 175924 279476 175976
rect 431960 175924 432012 175976
rect 273628 174768 273680 174820
rect 367100 174768 367152 174820
rect 273720 174700 273772 174752
rect 371240 174700 371292 174752
rect 275100 174632 275152 174684
rect 378140 174632 378192 174684
rect 280620 174564 280672 174616
rect 454040 174564 454092 174616
rect 287336 174496 287388 174548
rect 539692 174496 539744 174548
rect 292120 173476 292172 173528
rect 404360 173476 404412 173528
rect 285864 173408 285916 173460
rect 520280 173408 520332 173460
rect 285956 173340 286008 173392
rect 527180 173340 527232 173392
rect 287244 173272 287296 173324
rect 540980 173272 541032 173324
rect 288716 173204 288768 173256
rect 563060 173204 563112 173256
rect 289912 173136 289964 173188
rect 576860 173136 576912 173188
rect 291936 172320 291988 172372
rect 393320 172320 393372 172372
rect 292028 172252 292080 172304
rect 397460 172252 397512 172304
rect 295984 172184 296036 172236
rect 456892 172184 456944 172236
rect 283472 172116 283524 172168
rect 484400 172116 484452 172168
rect 283288 172048 283340 172100
rect 488540 172048 488592 172100
rect 283196 171980 283248 172032
rect 490012 171980 490064 172032
rect 283380 171912 283432 171964
rect 492680 171912 492732 171964
rect 284668 171844 284720 171896
rect 506480 171844 506532 171896
rect 284760 171776 284812 171828
rect 513380 171776 513432 171828
rect 276756 170756 276808 170808
rect 364340 170756 364392 170808
rect 293408 170688 293460 170740
rect 422300 170688 422352 170740
rect 279148 170620 279200 170672
rect 432052 170620 432104 170672
rect 279240 170552 279292 170604
rect 434720 170552 434772 170604
rect 279332 170484 279384 170536
rect 441620 170484 441672 170536
rect 282000 170416 282052 170468
rect 473360 170416 473412 170468
rect 282092 170348 282144 170400
rect 476120 170348 476172 170400
rect 273904 169192 273956 169244
rect 349344 169192 349396 169244
rect 280528 169124 280580 169176
rect 462320 169124 462372 169176
rect 281908 169056 281960 169108
rect 469220 169056 469272 169108
rect 283104 168988 283156 169040
rect 485780 168988 485832 169040
rect 278872 168104 278924 168156
rect 433340 168104 433392 168156
rect 279056 168036 279108 168088
rect 437480 168036 437532 168088
rect 278964 167968 279016 168020
rect 440240 167968 440292 168020
rect 280344 167900 280396 167952
rect 455420 167900 455472 167952
rect 280436 167832 280488 167884
rect 458180 167832 458232 167884
rect 280252 167764 280304 167816
rect 460940 167764 460992 167816
rect 281816 167696 281868 167748
rect 478880 167696 478932 167748
rect 289820 167628 289872 167680
rect 582380 167628 582432 167680
rect 407764 166948 407816 167000
rect 580172 166948 580224 167000
rect 277584 166608 277636 166660
rect 412640 166608 412692 166660
rect 293316 166540 293368 166592
rect 429200 166540 429252 166592
rect 277400 166472 277452 166524
rect 415492 166472 415544 166524
rect 277492 166404 277544 166456
rect 419540 166404 419592 166456
rect 278780 166336 278832 166388
rect 440332 166336 440384 166388
rect 291844 166268 291896 166320
rect 554780 166268 554832 166320
rect 274732 165248 274784 165300
rect 382372 165248 382424 165300
rect 274824 165180 274876 165232
rect 383660 165180 383712 165232
rect 274916 165112 274968 165164
rect 387800 165112 387852 165164
rect 275008 165044 275060 165096
rect 390652 165044 390704 165096
rect 276204 164976 276256 165028
rect 400220 164976 400272 165028
rect 276112 164908 276164 164960
rect 401600 164908 401652 164960
rect 276020 164840 276072 164892
rect 405740 164840 405792 164892
rect 3332 164160 3384 164212
rect 234804 164160 234856 164212
rect 273444 163888 273496 163940
rect 362960 163888 363012 163940
rect 273352 163820 273404 163872
rect 365812 163820 365864 163872
rect 273536 163752 273588 163804
rect 369860 163752 369912 163804
rect 256424 163684 256476 163736
rect 357440 163684 357492 163736
rect 274640 163616 274692 163668
rect 380900 163616 380952 163668
rect 311164 163548 311216 163600
rect 581092 163548 581144 163600
rect 234804 163480 234856 163532
rect 235540 163480 235592 163532
rect 272616 163480 272668 163532
rect 288624 163480 288676 163532
rect 558920 163480 558972 163532
rect 276664 162256 276716 162308
rect 372620 162256 372672 162308
rect 284576 162188 284628 162240
rect 506572 162188 506624 162240
rect 272616 162120 272668 162172
rect 285772 162120 285824 162172
rect 288532 162120 288584 162172
rect 564532 162120 564584 162172
rect 242624 161372 242676 161424
rect 267004 161372 267056 161424
rect 245476 161304 245528 161356
rect 269948 161304 270000 161356
rect 259552 161236 259604 161288
rect 299480 161236 299532 161288
rect 242716 161168 242768 161220
rect 267188 161168 267240 161220
rect 272524 161168 272576 161220
rect 347964 161168 348016 161220
rect 244004 161100 244056 161152
rect 268568 161100 268620 161152
rect 271236 161100 271288 161152
rect 348240 161100 348292 161152
rect 242072 161032 242124 161084
rect 267096 161032 267148 161084
rect 272432 161032 272484 161084
rect 350540 161032 350592 161084
rect 241336 160964 241388 161016
rect 268016 160964 268068 161016
rect 281448 160964 281500 161016
rect 448612 160964 448664 161016
rect 239956 160896 240008 160948
rect 268292 160896 268344 160948
rect 281724 160896 281776 160948
rect 477500 160896 477552 160948
rect 239680 160828 239732 160880
rect 268108 160828 268160 160880
rect 287152 160828 287204 160880
rect 543740 160828 543792 160880
rect 239772 160760 239824 160812
rect 268476 160760 268528 160812
rect 287060 160760 287112 160812
rect 547972 160760 548024 160812
rect 44180 160692 44232 160744
rect 247684 160692 247736 160744
rect 250996 160692 251048 160744
rect 268384 160692 268436 160744
rect 288440 160692 288492 160744
rect 561680 160692 561732 160744
rect 242808 160624 242860 160676
rect 265440 160624 265492 160676
rect 246856 160556 246908 160608
rect 268200 160556 268252 160608
rect 248696 160488 248748 160540
rect 264152 160488 264204 160540
rect 251640 159808 251692 159860
rect 263968 159808 264020 159860
rect 247592 159740 247644 159792
rect 264060 159740 264112 159792
rect 244464 159672 244516 159724
rect 263876 159672 263928 159724
rect 230480 159604 230532 159656
rect 262496 159604 262548 159656
rect 223580 159536 223632 159588
rect 262404 159536 262456 159588
rect 300400 159536 300452 159588
rect 327632 159536 327684 159588
rect 382924 159536 382976 159588
rect 465172 159536 465224 159588
rect 222200 159468 222252 159520
rect 262588 159468 262640 159520
rect 281632 159468 281684 159520
rect 470600 159468 470652 159520
rect 212540 159400 212592 159452
rect 261300 159400 261352 159452
rect 286692 159400 286744 159452
rect 525800 159400 525852 159452
rect 176752 159332 176804 159384
rect 258356 159332 258408 159384
rect 285864 159332 285916 159384
rect 529940 159332 529992 159384
rect 255228 158652 255280 158704
rect 269396 158652 269448 158704
rect 272892 158652 272944 158704
rect 300860 158652 300912 158704
rect 301504 158652 301556 158704
rect 345572 158652 345624 158704
rect 249708 158584 249760 158636
rect 265348 158584 265400 158636
rect 272064 158584 272116 158636
rect 346952 158584 347004 158636
rect 251088 158516 251140 158568
rect 266820 158516 266872 158568
rect 271144 158516 271196 158568
rect 348056 158516 348108 158568
rect 249616 158448 249668 158500
rect 267924 158448 267976 158500
rect 272248 158448 272300 158500
rect 349712 158448 349764 158500
rect 246672 158380 246724 158432
rect 266728 158380 266780 158432
rect 270960 158380 271012 158432
rect 349528 158380 349580 158432
rect 246764 158312 246816 158364
rect 242992 158244 243044 158296
rect 263784 158244 263836 158296
rect 264520 158312 264572 158364
rect 265624 158312 265676 158364
rect 271052 158312 271104 158364
rect 349804 158312 349856 158364
rect 266912 158244 266964 158296
rect 269488 158244 269540 158296
rect 349620 158244 349672 158296
rect 219440 158176 219492 158228
rect 262864 158176 262916 158228
rect 272156 158176 272208 158228
rect 353300 158176 353352 158228
rect 208400 158108 208452 158160
rect 261208 158108 261260 158160
rect 271972 158108 272024 158160
rect 357532 158108 357584 158160
rect 204260 158040 204312 158092
rect 261116 158040 261168 158092
rect 284484 158040 284536 158092
rect 187700 157972 187752 158024
rect 259828 157972 259880 158024
rect 259920 157972 259972 158024
rect 260564 157972 260616 158024
rect 281264 157972 281316 158024
rect 287704 157972 287756 158024
rect 293224 158040 293276 158092
rect 411260 158040 411312 158092
rect 505100 157972 505152 158024
rect 253848 157904 253900 157956
rect 266636 157904 266688 157956
rect 301688 157904 301740 157956
rect 331496 157904 331548 157956
rect 337384 157904 337436 157956
rect 339868 157904 339920 157956
rect 300308 157836 300360 157888
rect 319260 157836 319312 157888
rect 256792 157768 256844 157820
rect 261484 157768 261536 157820
rect 301596 157768 301648 157820
rect 314752 157768 314804 157820
rect 259828 157428 259880 157480
rect 265256 157428 265308 157480
rect 3608 157360 3660 157412
rect 293960 157360 294012 157412
rect 250444 156884 250496 156936
rect 264244 157020 264296 157072
rect 240140 156816 240192 156868
rect 264336 156952 264388 157004
rect 300124 156952 300176 157004
rect 345020 156952 345072 157004
rect 300216 156884 300268 156936
rect 345756 156884 345808 156936
rect 231860 156748 231912 156800
rect 262680 156816 262732 156868
rect 273260 156816 273312 156868
rect 360200 156816 360252 156868
rect 213920 156680 213972 156732
rect 261024 156748 261076 156800
rect 281540 156748 281592 156800
rect 473452 156748 473504 156800
rect 259644 156680 259696 156732
rect 265164 156680 265216 156732
rect 283012 156680 283064 156732
rect 495440 156680 495492 156732
rect 205640 156612 205692 156664
rect 259736 156612 259788 156664
rect 260748 156612 260800 156664
rect 285312 156612 285364 156664
rect 502340 156612 502392 156664
rect 261668 156544 261720 156596
rect 259920 156000 259972 156052
rect 260380 156000 260432 156052
rect 259276 155864 259328 155916
rect 265532 155864 265584 155916
rect 259092 155796 259144 155848
rect 266544 155796 266596 155848
rect 270868 155796 270920 155848
rect 259184 155728 259236 155780
rect 267556 155728 267608 155780
rect 270776 155728 270828 155780
rect 260288 155660 260340 155712
rect 261576 155660 261628 155712
rect 270684 155660 270736 155712
rect 271880 155660 271932 155712
rect 257712 155592 257764 155644
rect 267832 155592 267884 155644
rect 269120 155592 269172 155644
rect 257528 155524 257580 155576
rect 268660 155524 268712 155576
rect 253756 155456 253808 155508
rect 265808 155456 265860 155508
rect 197360 155388 197412 155440
rect 260012 155388 260064 155440
rect 260472 155388 260524 155440
rect 270592 155388 270644 155440
rect 194600 155320 194652 155372
rect 259460 155320 259512 155372
rect 193312 155252 193364 155304
rect 190460 155184 190512 155236
rect 259920 155184 259972 155236
rect 271696 155388 271748 155440
rect 344192 155524 344244 155576
rect 344376 155456 344428 155508
rect 271880 155388 271932 155440
rect 344468 155388 344520 155440
rect 344560 155320 344612 155372
rect 347136 155252 347188 155304
rect 347228 155184 347280 155236
rect 30380 153824 30432 153876
rect 247500 153824 247552 153876
rect 233976 153144 234028 153196
rect 256700 153144 256752 153196
rect 3332 150356 3384 150408
rect 94504 150356 94556 150408
rect 234160 144848 234212 144900
rect 256700 144848 256752 144900
rect 257252 142060 257304 142112
rect 257804 142060 257856 142112
rect 577688 139340 577740 139392
rect 579620 139340 579672 139392
rect 3056 137912 3108 137964
rect 235264 137912 235316 137964
rect 234252 135192 234304 135244
rect 256792 135192 256844 135244
rect 232504 131044 232556 131096
rect 256792 131044 256844 131096
rect 344284 130364 344336 130416
rect 345020 130364 345072 130416
rect 234804 126896 234856 126948
rect 235632 126896 235684 126948
rect 256792 126896 256844 126948
rect 347044 126896 347096 126948
rect 579712 126896 579764 126948
rect 90456 126216 90508 126268
rect 234804 126216 234856 126268
rect 235724 122748 235776 122800
rect 256792 122748 256844 122800
rect 234344 113092 234396 113144
rect 256792 113092 256844 113144
rect 234528 104796 234580 104848
rect 256792 104796 256844 104848
rect 577596 100648 577648 100700
rect 579620 100648 579672 100700
rect 259736 100444 259788 100496
rect 263692 100444 263744 100496
rect 256516 100036 256568 100088
rect 260840 100036 260892 100088
rect 246948 99968 247000 100020
rect 262220 99968 262272 100020
rect 257988 97928 258040 97980
rect 267740 97928 267792 97980
rect 334716 97928 334768 97980
rect 349896 97928 349948 97980
rect 245108 97860 245160 97912
rect 297364 97860 297416 97912
rect 317972 97860 318024 97912
rect 349252 97860 349304 97912
rect 259000 97792 259052 97844
rect 301228 97792 301280 97844
rect 339224 97792 339276 97844
rect 347872 97792 347924 97844
rect 257896 97724 257948 97776
rect 276112 97724 276164 97776
rect 322480 97724 322532 97776
rect 347780 97724 347832 97776
rect 259552 97656 259604 97708
rect 284484 97656 284536 97708
rect 326344 97656 326396 97708
rect 348332 97656 348384 97708
rect 257344 97588 257396 97640
rect 280620 97588 280672 97640
rect 309600 97588 309652 97640
rect 344652 97588 344704 97640
rect 234436 97520 234488 97572
rect 292856 97520 292908 97572
rect 314108 97520 314160 97572
rect 344008 97520 344060 97572
rect 235816 97452 235868 97504
rect 263876 97452 263928 97504
rect 99380 89020 99432 89072
rect 243820 89020 243872 89072
rect 92480 88952 92532 89004
rect 243912 88952 243964 89004
rect 3332 85484 3384 85536
rect 90364 85484 90416 85536
rect 86960 82084 87012 82136
rect 251548 82084 251600 82136
rect 3332 71680 3384 71732
rect 235908 71680 235960 71732
rect 305000 71680 305052 71732
rect 3332 59304 3384 59356
rect 231124 59304 231176 59356
rect 3516 33056 3568 33108
rect 90456 33056 90508 33108
rect 142160 21360 142212 21412
rect 255596 21360 255648 21412
rect 3516 20612 3568 20664
rect 174544 20612 174596 20664
rect 577504 20612 577556 20664
rect 579712 20612 579764 20664
rect 120632 14560 120684 14612
rect 254308 14560 254360 14612
rect 110512 14492 110564 14544
rect 253020 14492 253072 14544
rect 102232 14424 102284 14476
rect 252928 14424 252980 14476
rect 124680 13200 124732 13252
rect 245016 13200 245068 13252
rect 122288 13132 122340 13184
rect 254216 13132 254268 13184
rect 13544 13064 13596 13116
rect 246028 13064 246080 13116
rect 127624 12248 127676 12300
rect 250352 12248 250404 12300
rect 117320 12180 117372 12232
rect 254124 12180 254176 12232
rect 108120 12112 108172 12164
rect 252652 12112 252704 12164
rect 104072 12044 104124 12096
rect 252836 12044 252888 12096
rect 100760 11976 100812 12028
rect 252744 11976 252796 12028
rect 89904 11908 89956 11960
rect 251456 11908 251508 11960
rect 5264 11840 5316 11892
rect 178868 11840 178920 11892
rect 347964 11840 348016 11892
rect 73344 11772 73396 11824
rect 250260 11772 250312 11824
rect 33600 11704 33652 11756
rect 247408 11704 247460 11756
rect 160100 11636 160152 11688
rect 161296 11636 161348 11688
rect 184940 11636 184992 11688
rect 186136 11636 186188 11688
rect 201500 11636 201552 11688
rect 202696 11636 202748 11688
rect 234620 11636 234672 11688
rect 235816 11636 235868 11688
rect 348056 11636 348108 11688
rect 181444 10684 181496 10736
rect 251364 10684 251416 10736
rect 114008 10616 114060 10668
rect 242532 10616 242584 10668
rect 42800 10548 42852 10600
rect 200764 10548 200816 10600
rect 20168 10480 20220 10532
rect 182824 10480 182876 10532
rect 221464 10480 221516 10532
rect 247224 10480 247276 10532
rect 69112 10412 69164 10464
rect 250168 10412 250220 10464
rect 36728 10344 36780 10396
rect 247316 10344 247368 10396
rect 11888 10276 11940 10328
rect 245936 10276 245988 10328
rect 239680 9596 239732 9648
rect 291384 9596 291436 9648
rect 196072 9528 196124 9580
rect 250076 9528 250128 9580
rect 239772 9460 239824 9512
rect 294880 9460 294932 9512
rect 239956 9392 240008 9444
rect 298468 9392 298520 9444
rect 241336 9324 241388 9376
rect 301964 9324 302016 9376
rect 239588 9256 239640 9308
rect 305552 9256 305604 9308
rect 241244 9188 241296 9240
rect 309048 9188 309100 9240
rect 239864 9120 239916 9172
rect 312636 9120 312688 9172
rect 138848 9052 138900 9104
rect 251824 9052 251876 9104
rect 106924 8984 106976 9036
rect 242440 8984 242492 9036
rect 244004 8984 244056 9036
rect 287796 8984 287848 9036
rect 35992 8916 36044 8968
rect 196624 8916 196676 8968
rect 241152 8916 241204 8968
rect 316224 8916 316276 8968
rect 240048 8848 240100 8900
rect 284300 8848 284352 8900
rect 242072 8780 242124 8832
rect 280712 8780 280764 8832
rect 242624 8712 242676 8764
rect 277124 8712 277176 8764
rect 170772 8032 170824 8084
rect 258724 8032 258776 8084
rect 143540 7964 143592 8016
rect 255504 7964 255556 8016
rect 103336 7896 103388 7948
rect 253664 7896 253716 7948
rect 85672 7828 85724 7880
rect 243728 7828 243780 7880
rect 28908 7760 28960 7812
rect 188344 7760 188396 7812
rect 199108 7760 199160 7812
rect 254584 7760 254636 7812
rect 11152 7692 11204 7744
rect 178684 7692 178736 7744
rect 180248 7692 180300 7744
rect 258264 7692 258316 7744
rect 83280 7624 83332 7676
rect 252100 7624 252152 7676
rect 51356 7556 51408 7608
rect 249524 7556 249576 7608
rect 246764 6808 246816 6860
rect 279516 6808 279568 6860
rect 344928 6808 344980 6860
rect 580172 6808 580224 6860
rect 246672 6740 246724 6792
rect 283104 6740 283156 6792
rect 248328 6672 248380 6724
rect 286600 6672 286652 6724
rect 244096 6604 244148 6656
rect 293684 6604 293736 6656
rect 246856 6536 246908 6588
rect 300768 6536 300820 6588
rect 248236 6468 248288 6520
rect 304356 6468 304408 6520
rect 245476 6400 245528 6452
rect 307944 6400 307996 6452
rect 173164 6332 173216 6384
rect 258540 6332 258592 6384
rect 78588 6264 78640 6316
rect 249156 6264 249208 6316
rect 249616 6264 249668 6316
rect 290188 6264 290240 6316
rect 72608 6196 72660 6248
rect 249984 6196 250036 6248
rect 250996 6196 251048 6248
rect 297272 6196 297324 6248
rect 337476 6196 337528 6248
rect 348240 6196 348292 6248
rect 19432 6128 19484 6180
rect 242348 6128 242400 6180
rect 245568 6128 245620 6180
rect 311440 6128 311492 6180
rect 333888 6128 333940 6180
rect 349804 6128 349856 6180
rect 242716 6060 242768 6112
rect 273628 6060 273680 6112
rect 241428 5992 241480 6044
rect 270040 5992 270092 6044
rect 242808 5924 242860 5976
rect 266544 5924 266596 5976
rect 197360 5108 197412 5160
rect 255780 5108 255832 5160
rect 175924 5040 175976 5092
rect 244280 5040 244332 5092
rect 64328 4972 64380 5024
rect 250812 4972 250864 5024
rect 57244 4904 57296 4956
rect 248972 4904 249024 4956
rect 14740 4836 14792 4888
rect 246212 4836 246264 4888
rect 1676 4768 1728 4820
rect 244372 4768 244424 4820
rect 253848 4088 253900 4140
rect 272432 4088 272484 4140
rect 329196 4088 329248 4140
rect 347228 4088 347280 4140
rect 249708 4020 249760 4072
rect 268844 4020 268896 4072
rect 328000 4020 328052 4072
rect 346676 4020 346728 4072
rect 259184 3952 259236 4004
rect 281908 3952 281960 4004
rect 325608 3952 325660 4004
rect 344376 3952 344428 4004
rect 128176 3884 128228 3936
rect 182916 3884 182968 3936
rect 251088 3884 251140 3936
rect 276020 3884 276072 3936
rect 324412 3884 324464 3936
rect 346768 3884 346820 3936
rect 141240 3816 141292 3868
rect 197360 3816 197412 3868
rect 203892 3816 203944 3868
rect 243544 3816 243596 3868
rect 257620 3816 257672 3868
rect 285404 3816 285456 3868
rect 322112 3816 322164 3868
rect 345848 3816 345900 3868
rect 70308 3748 70360 3800
rect 127624 3748 127676 3800
rect 175464 3748 175516 3800
rect 249064 3748 249116 3800
rect 257712 3748 257764 3800
rect 288992 3748 289044 3800
rect 320916 3748 320968 3800
rect 343916 3748 343968 3800
rect 86868 3680 86920 3732
rect 181444 3680 181496 3732
rect 196808 3680 196860 3732
rect 243636 3680 243688 3732
rect 244188 3680 244240 3732
rect 278320 3680 278372 3732
rect 326804 3680 326856 3732
rect 349528 3680 349580 3732
rect 65524 3612 65576 3664
rect 196072 3612 196124 3664
rect 200304 3612 200356 3664
rect 242164 3612 242216 3664
rect 259368 3612 259420 3664
rect 296076 3612 296128 3664
rect 323308 3612 323360 3664
rect 348148 3612 348200 3664
rect 2872 3544 2924 3596
rect 175924 3544 175976 3596
rect 179052 3544 179104 3596
rect 233884 3544 233936 3596
rect 244924 3544 244976 3596
rect 256608 3544 256660 3596
rect 292580 3544 292632 3596
rect 318524 3544 318576 3596
rect 344652 3544 344704 3596
rect 30104 3476 30156 3528
rect 221464 3476 221516 3528
rect 226340 3476 226392 3528
rect 227536 3476 227588 3528
rect 227628 3476 227680 3528
rect 242256 3476 242308 3528
rect 15936 3408 15988 3460
rect 254676 3476 254728 3528
rect 256056 3476 256108 3528
rect 257528 3476 257580 3528
rect 299664 3476 299716 3528
rect 319720 3476 319772 3528
rect 349620 3544 349672 3596
rect 365812 3476 365864 3528
rect 367008 3476 367060 3528
rect 374092 3476 374144 3528
rect 375288 3476 375340 3528
rect 382372 3476 382424 3528
rect 383568 3476 383620 3528
rect 390652 3476 390704 3528
rect 391848 3476 391900 3528
rect 407212 3476 407264 3528
rect 408408 3476 408460 3528
rect 415492 3476 415544 3528
rect 416688 3476 416740 3528
rect 423772 3476 423824 3528
rect 424968 3476 425020 3528
rect 432052 3476 432104 3528
rect 433248 3476 433300 3528
rect 448612 3476 448664 3528
rect 449808 3476 449860 3528
rect 456892 3476 456944 3528
rect 458088 3476 458140 3528
rect 465080 3476 465132 3528
rect 465908 3476 465960 3528
rect 489920 3476 489972 3528
rect 490748 3476 490800 3528
rect 498200 3476 498252 3528
rect 499028 3476 499080 3528
rect 514760 3476 514812 3528
rect 515588 3476 515640 3528
rect 523040 3476 523092 3528
rect 523868 3476 523920 3528
rect 539600 3476 539652 3528
rect 540428 3476 540480 3528
rect 547880 3476 547932 3528
rect 548708 3476 548760 3528
rect 581000 3476 581052 3528
rect 581828 3476 581880 3528
rect 246396 3408 246448 3460
rect 254584 3408 254636 3460
rect 257436 3408 257488 3460
rect 303160 3408 303212 3460
rect 315028 3408 315080 3460
rect 346400 3408 346452 3460
rect 356704 3408 356756 3460
rect 579804 3408 579856 3460
rect 44180 3340 44232 3392
rect 45100 3340 45152 3392
rect 259092 3340 259144 3392
rect 271236 3340 271288 3392
rect 330392 3340 330444 3392
rect 347872 3340 347924 3392
rect 253756 3272 253808 3324
rect 265348 3272 265400 3324
rect 331588 3272 331640 3324
rect 346584 3272 346636 3324
rect 259276 3204 259328 3256
rect 267740 3204 267792 3256
rect 332692 3204 332744 3256
rect 346860 3204 346912 3256
rect 252376 3136 252428 3188
rect 255964 3136 256016 3188
rect 226340 2796 226392 2848
rect 227628 2796 227680 2848
rect 357440 2184 357492 2236
rect 358728 2184 358780 2236
rect 398840 2184 398892 2236
rect 400128 2184 400180 2236
rect 440240 2184 440292 2236
rect 441528 2184 441580 2236
<< metal2 >>
rect 6932 703582 7972 703610
rect 3422 684312 3478 684321
rect 3422 684247 3478 684256
rect 3436 683262 3464 684247
rect 3424 683256 3476 683262
rect 3424 683198 3476 683204
rect 3422 671256 3478 671265
rect 3422 671191 3478 671200
rect 3436 670818 3464 671191
rect 3424 670812 3476 670818
rect 3424 670754 3476 670760
rect 3422 658200 3478 658209
rect 3422 658135 3478 658144
rect 3436 656946 3464 658135
rect 3424 656940 3476 656946
rect 3424 656882 3476 656888
rect 3424 632120 3476 632126
rect 3422 632088 3424 632097
rect 3476 632088 3478 632097
rect 3422 632023 3478 632032
rect 2778 619168 2834 619177
rect 2778 619103 2780 619112
rect 2832 619103 2834 619112
rect 4804 619132 4856 619138
rect 2780 619074 2832 619080
rect 4804 619074 4856 619080
rect 3238 606112 3294 606121
rect 3238 606047 3294 606056
rect 3252 605878 3280 606047
rect 3240 605872 3292 605878
rect 3240 605814 3292 605820
rect 3422 580000 3478 580009
rect 3422 579935 3478 579944
rect 2778 566944 2834 566953
rect 2778 566879 2834 566888
rect 2792 566098 2820 566879
rect 2780 566092 2832 566098
rect 2780 566034 2832 566040
rect 2778 553888 2834 553897
rect 2778 553823 2834 553832
rect 2792 553722 2820 553823
rect 2780 553716 2832 553722
rect 2780 553658 2832 553664
rect 3330 501800 3386 501809
rect 3330 501735 3386 501744
rect 3344 501362 3372 501735
rect 3332 501356 3384 501362
rect 3332 501298 3384 501304
rect 3330 475688 3386 475697
rect 3330 475623 3386 475632
rect 3344 474774 3372 475623
rect 3332 474768 3384 474774
rect 3332 474710 3384 474716
rect 3330 462632 3386 462641
rect 3330 462567 3386 462576
rect 3344 462398 3372 462567
rect 3332 462392 3384 462398
rect 3332 462334 3384 462340
rect 3330 449576 3386 449585
rect 3330 449511 3386 449520
rect 3344 448594 3372 449511
rect 3332 448588 3384 448594
rect 3332 448530 3384 448536
rect 3146 423600 3202 423609
rect 3146 423535 3202 423544
rect 3160 422346 3188 423535
rect 3148 422340 3200 422346
rect 3148 422282 3200 422288
rect 3146 410544 3202 410553
rect 3146 410479 3202 410488
rect 3160 409902 3188 410479
rect 3148 409896 3200 409902
rect 3148 409838 3200 409844
rect 3332 397520 3384 397526
rect 3330 397488 3332 397497
rect 3384 397488 3386 397497
rect 3330 397423 3386 397432
rect 3436 387258 3464 579935
rect 3514 527912 3570 527921
rect 3514 527847 3570 527856
rect 3528 388482 3556 527847
rect 3606 514856 3662 514865
rect 3606 514791 3662 514800
rect 3620 393990 3648 514791
rect 3608 393984 3660 393990
rect 4816 393961 4844 619074
rect 4896 566092 4948 566098
rect 4896 566034 4948 566040
rect 3608 393926 3660 393932
rect 4802 393952 4858 393961
rect 4802 393887 4858 393896
rect 4908 388550 4936 566034
rect 4988 553716 5040 553722
rect 4988 553658 5040 553664
rect 5000 391270 5028 553658
rect 6932 391338 6960 703582
rect 7944 703474 7972 703582
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40052 703582 40356 703610
rect 8128 703474 8156 703520
rect 7944 703446 8156 703474
rect 24320 700330 24348 703520
rect 24308 700324 24360 700330
rect 24308 700266 24360 700272
rect 7564 501356 7616 501362
rect 7564 501298 7616 501304
rect 7576 392766 7604 501298
rect 7564 392760 7616 392766
rect 7564 392702 7616 392708
rect 6920 391332 6972 391338
rect 6920 391274 6972 391280
rect 4988 391264 5040 391270
rect 4988 391206 5040 391212
rect 40052 388686 40080 703582
rect 40328 703474 40356 703582
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 104912 703582 105308 703610
rect 40512 703474 40540 703520
rect 40328 703446 40540 703474
rect 72988 703050 73016 703520
rect 71780 703044 71832 703050
rect 71780 702986 71832 702992
rect 72976 703044 73028 703050
rect 72976 702986 73028 702992
rect 71792 389978 71820 702986
rect 89180 700398 89208 703520
rect 89168 700392 89220 700398
rect 89168 700334 89220 700340
rect 104912 590034 104940 703582
rect 105280 703474 105308 703582
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 136652 703582 137692 703610
rect 105464 703474 105492 703520
rect 105280 703446 105492 703474
rect 136652 590102 136680 703582
rect 137664 703474 137692 703582
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 234632 703582 235028 703610
rect 137848 703474 137876 703520
rect 137664 703446 137876 703474
rect 154132 700466 154160 703520
rect 170324 700534 170352 703520
rect 202800 703050 202828 703520
rect 201500 703044 201552 703050
rect 201500 702986 201552 702992
rect 202788 703044 202840 703050
rect 202788 702986 202840 702992
rect 170312 700528 170364 700534
rect 170312 700470 170364 700476
rect 192484 700528 192536 700534
rect 192484 700470 192536 700476
rect 154120 700460 154172 700466
rect 154120 700402 154172 700408
rect 136640 590096 136692 590102
rect 136640 590038 136692 590044
rect 104900 590028 104952 590034
rect 104900 589970 104952 589976
rect 97814 537024 97870 537033
rect 97814 536959 97870 536968
rect 97630 510232 97686 510241
rect 97630 510167 97686 510176
rect 97538 508328 97594 508337
rect 97538 508263 97594 508272
rect 97552 426426 97580 508263
rect 97540 426420 97592 426426
rect 97540 426362 97592 426368
rect 97644 397458 97672 510167
rect 97722 508600 97778 508609
rect 97722 508535 97778 508544
rect 97632 397452 97684 397458
rect 97632 397394 97684 397400
rect 71780 389972 71832 389978
rect 71780 389914 71832 389920
rect 40040 388680 40092 388686
rect 40040 388622 40092 388628
rect 4896 388544 4948 388550
rect 4896 388486 4948 388492
rect 3516 388476 3568 388482
rect 3516 388418 3568 388424
rect 3424 387252 3476 387258
rect 3424 387194 3476 387200
rect 97736 386374 97764 508535
rect 97828 398138 97856 536959
rect 97906 535936 97962 535945
rect 97906 535871 97962 535880
rect 97816 398132 97868 398138
rect 97816 398074 97868 398080
rect 97724 386368 97776 386374
rect 97724 386310 97776 386316
rect 97920 385694 97948 535871
rect 99194 534304 99250 534313
rect 99194 534239 99250 534248
rect 99102 533216 99158 533225
rect 99102 533151 99158 533160
rect 99010 530224 99066 530233
rect 99010 530159 99066 530168
rect 98918 528592 98974 528601
rect 98918 528527 98974 528536
rect 98932 396030 98960 528527
rect 98920 396024 98972 396030
rect 98920 395966 98972 395972
rect 99024 395962 99052 530159
rect 99116 397390 99144 533151
rect 99104 397384 99156 397390
rect 99104 397326 99156 397332
rect 99208 396778 99236 534239
rect 99286 531584 99342 531593
rect 99286 531519 99342 531528
rect 99196 396772 99248 396778
rect 99196 396714 99248 396720
rect 99012 395956 99064 395962
rect 99012 395898 99064 395904
rect 99300 385762 99328 531519
rect 114466 498128 114522 498137
rect 114466 498063 114522 498072
rect 119342 498128 119398 498137
rect 119342 498063 119398 498072
rect 123390 498128 123446 498137
rect 125230 498128 125286 498137
rect 123390 498063 123392 498072
rect 113086 496904 113142 496913
rect 113086 496839 113142 496848
rect 113100 394058 113128 496839
rect 114480 395350 114508 498063
rect 119356 497078 119384 498063
rect 123444 498063 123446 498072
rect 124864 498092 124916 498098
rect 123392 498034 123444 498040
rect 125230 498063 125286 498072
rect 126794 498128 126850 498137
rect 126794 498063 126850 498072
rect 151726 498128 151782 498137
rect 151726 498063 151782 498072
rect 124864 498034 124916 498040
rect 121366 497448 121422 497457
rect 121366 497383 121422 497392
rect 119344 497072 119396 497078
rect 119344 497014 119396 497020
rect 115478 496904 115534 496913
rect 118606 496904 118662 496913
rect 115478 496839 115480 496848
rect 115532 496839 115534 496848
rect 116584 496868 116636 496874
rect 115480 496810 115532 496816
rect 118606 496839 118662 496848
rect 121274 496904 121330 496913
rect 121274 496839 121330 496848
rect 116584 496810 116636 496816
rect 116596 395418 116624 496810
rect 118620 399566 118648 496839
rect 121288 400994 121316 496839
rect 121276 400988 121328 400994
rect 121276 400930 121328 400936
rect 118608 399560 118660 399566
rect 118608 399502 118660 399508
rect 121380 399498 121408 497383
rect 122746 496904 122802 496913
rect 122746 496839 122802 496848
rect 122760 400926 122788 496839
rect 124876 401062 124904 498034
rect 125244 496942 125272 498063
rect 126808 497010 126836 498063
rect 126796 497004 126848 497010
rect 126796 496946 126848 496952
rect 125232 496936 125284 496942
rect 125232 496878 125284 496884
rect 125506 496904 125562 496913
rect 125506 496839 125562 496848
rect 131026 496904 131082 496913
rect 131026 496839 131082 496848
rect 136546 496904 136602 496913
rect 136546 496839 136602 496848
rect 140686 496904 140742 496913
rect 140686 496839 140742 496848
rect 146206 496904 146262 496913
rect 146206 496839 146262 496848
rect 124864 401056 124916 401062
rect 124864 400998 124916 401004
rect 122748 400920 122800 400926
rect 122748 400862 122800 400868
rect 121368 399492 121420 399498
rect 121368 399434 121420 399440
rect 116584 395412 116636 395418
rect 116584 395354 116636 395360
rect 114468 395344 114520 395350
rect 114468 395286 114520 395292
rect 113088 394052 113140 394058
rect 113088 393994 113140 394000
rect 125520 385830 125548 496839
rect 131040 396846 131068 496839
rect 136560 398206 136588 496839
rect 140700 399634 140728 496839
rect 146220 414730 146248 496839
rect 151740 414798 151768 498063
rect 155866 496904 155922 496913
rect 155866 496839 155922 496848
rect 161386 496904 161442 496913
rect 161386 496839 161442 496848
rect 155880 414866 155908 496839
rect 155868 414860 155920 414866
rect 155868 414802 155920 414808
rect 151728 414792 151780 414798
rect 151728 414734 151780 414740
rect 146208 414724 146260 414730
rect 146208 414666 146260 414672
rect 161400 399702 161428 496839
rect 175924 462392 175976 462398
rect 175924 462334 175976 462340
rect 161388 399696 161440 399702
rect 161388 399638 161440 399644
rect 140688 399628 140740 399634
rect 140688 399570 140740 399576
rect 136548 398200 136600 398206
rect 136548 398142 136600 398148
rect 131028 396840 131080 396846
rect 131028 396782 131080 396788
rect 175936 385898 175964 462334
rect 192496 387394 192524 700470
rect 192576 700324 192628 700330
rect 192576 700266 192628 700272
rect 192588 392630 192616 700266
rect 192668 656940 192720 656946
rect 192668 656882 192720 656888
rect 192576 392624 192628 392630
rect 192576 392566 192628 392572
rect 192680 391610 192708 656882
rect 192668 391604 192720 391610
rect 192668 391546 192720 391552
rect 201512 388822 201540 702986
rect 218992 699718 219020 703520
rect 218980 699712 219032 699718
rect 218980 699654 219032 699660
rect 220084 699712 220136 699718
rect 220084 699654 220136 699660
rect 220096 392902 220124 699654
rect 234528 409896 234580 409902
rect 234528 409838 234580 409844
rect 233790 393952 233846 393961
rect 233790 393887 233846 393896
rect 233804 393417 233832 393887
rect 233790 393408 233846 393417
rect 233790 393343 233792 393352
rect 233844 393343 233846 393352
rect 233792 393314 233844 393320
rect 220084 392896 220136 392902
rect 220084 392838 220136 392844
rect 233976 392624 234028 392630
rect 233976 392566 234028 392572
rect 233988 392018 234016 392566
rect 233976 392012 234028 392018
rect 233976 391954 234028 391960
rect 233988 389450 234016 391954
rect 233988 389422 234108 389450
rect 201500 388816 201552 388822
rect 201500 388758 201552 388764
rect 192484 387388 192536 387394
rect 192484 387330 192536 387336
rect 175924 385892 175976 385898
rect 175924 385834 175976 385840
rect 125508 385824 125560 385830
rect 125508 385766 125560 385772
rect 99288 385756 99340 385762
rect 99288 385698 99340 385704
rect 97908 385688 97960 385694
rect 97908 385630 97960 385636
rect 174544 384668 174596 384674
rect 174544 384610 174596 384616
rect 3792 382968 3844 382974
rect 3792 382910 3844 382916
rect 3700 381608 3752 381614
rect 3700 381550 3752 381556
rect 3424 381540 3476 381546
rect 3424 381482 3476 381488
rect 3148 372564 3200 372570
rect 3148 372506 3200 372512
rect 3160 371385 3188 372506
rect 3146 371376 3202 371385
rect 3146 371311 3202 371320
rect 2964 346384 3016 346390
rect 2964 346326 3016 346332
rect 2976 345409 3004 346326
rect 2962 345400 3018 345409
rect 2962 345335 3018 345344
rect 20 323604 72 323610
rect 20 323546 72 323552
rect 32 16574 60 323546
rect 3148 320136 3200 320142
rect 3148 320078 3200 320084
rect 3160 319297 3188 320078
rect 3146 319288 3202 319297
rect 3146 319223 3202 319232
rect 3332 306332 3384 306338
rect 3332 306274 3384 306280
rect 3344 306241 3372 306274
rect 3330 306232 3386 306241
rect 3330 306167 3386 306176
rect 3240 293956 3292 293962
rect 3240 293898 3292 293904
rect 3252 293185 3280 293898
rect 3238 293176 3294 293185
rect 3238 293111 3294 293120
rect 3330 267200 3386 267209
rect 3330 267135 3386 267144
rect 3344 267034 3372 267135
rect 3332 267028 3384 267034
rect 3332 266970 3384 266976
rect 3332 255264 3384 255270
rect 3332 255206 3384 255212
rect 3344 254153 3372 255206
rect 3330 254144 3386 254153
rect 3330 254079 3386 254088
rect 3332 241460 3384 241466
rect 3332 241402 3384 241408
rect 3344 241097 3372 241402
rect 3330 241088 3386 241097
rect 3330 241023 3386 241032
rect 3330 214976 3386 214985
rect 3330 214911 3386 214920
rect 3344 214606 3372 214911
rect 3332 214600 3384 214606
rect 3332 214542 3384 214548
rect 2780 178696 2832 178702
rect 2780 178638 2832 178644
rect 2792 16574 2820 178638
rect 3332 164212 3384 164218
rect 3332 164154 3384 164160
rect 3344 162897 3372 164154
rect 3330 162888 3386 162897
rect 3330 162823 3386 162832
rect 3332 150408 3384 150414
rect 3332 150350 3384 150356
rect 3344 149841 3372 150350
rect 3330 149832 3386 149841
rect 3330 149767 3386 149776
rect 3056 137964 3108 137970
rect 3056 137906 3108 137912
rect 3068 136785 3096 137906
rect 3054 136776 3110 136785
rect 3054 136711 3110 136720
rect 3332 85536 3384 85542
rect 3332 85478 3384 85484
rect 3344 84697 3372 85478
rect 3330 84688 3386 84697
rect 3330 84623 3386 84632
rect 3332 71732 3384 71738
rect 3332 71674 3384 71680
rect 3344 71641 3372 71674
rect 3330 71632 3386 71641
rect 3330 71567 3386 71576
rect 3332 59356 3384 59362
rect 3332 59298 3384 59304
rect 3344 58585 3372 59298
rect 3330 58576 3386 58585
rect 3330 58511 3386 58520
rect 32 16546 152 16574
rect 2792 16546 3372 16574
rect 124 354 152 16546
rect 1676 4820 1728 4826
rect 1676 4762 1728 4768
rect 1688 480 1716 4762
rect 2872 3596 2924 3602
rect 2872 3538 2924 3544
rect 2884 480 2912 3538
rect 3344 490 3372 16546
rect 3436 6497 3464 381482
rect 3514 381168 3570 381177
rect 3514 381103 3570 381112
rect 3528 45529 3556 381103
rect 3608 381064 3660 381070
rect 3608 381006 3660 381012
rect 3620 188873 3648 381006
rect 3712 201929 3740 381550
rect 3804 358465 3832 382910
rect 90362 382664 90418 382673
rect 90362 382599 90418 382608
rect 3790 358456 3846 358465
rect 3790 358391 3846 358400
rect 81440 337340 81492 337346
rect 81440 337282 81492 337288
rect 26240 337272 26292 337278
rect 26240 337214 26292 337220
rect 24858 333296 24914 333305
rect 24858 333231 24914 333240
rect 9678 327720 9734 327729
rect 9678 327655 9734 327664
rect 6918 326360 6974 326369
rect 6918 326295 6974 326304
rect 3698 201920 3754 201929
rect 3698 201855 3754 201864
rect 3606 188864 3662 188873
rect 3606 188799 3662 188808
rect 3608 157412 3660 157418
rect 3608 157354 3660 157360
rect 3620 110673 3648 157354
rect 3606 110664 3662 110673
rect 3606 110599 3662 110608
rect 3514 45520 3570 45529
rect 3514 45455 3570 45464
rect 3516 33108 3568 33114
rect 3516 33050 3568 33056
rect 3528 32473 3556 33050
rect 3514 32464 3570 32473
rect 3514 32399 3570 32408
rect 3516 20664 3568 20670
rect 3516 20606 3568 20612
rect 3528 19417 3556 20606
rect 3514 19408 3570 19417
rect 3514 19343 3570 19352
rect 6932 16574 6960 326295
rect 6932 16546 7696 16574
rect 5264 11892 5316 11898
rect 5264 11834 5316 11840
rect 3422 6488 3478 6497
rect 3422 6423 3478 6432
rect 542 354 654 480
rect 124 326 654 354
rect 542 -960 654 326
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 3344 462 3740 490
rect 5276 480 5304 11834
rect 6458 4856 6514 4865
rect 6458 4791 6514 4800
rect 6472 480 6500 4791
rect 7668 480 7696 16546
rect 8758 13016 8814 13025
rect 8758 12951 8814 12960
rect 8772 480 8800 12951
rect 3712 354 3740 462
rect 4038 354 4150 480
rect 3712 326 4150 354
rect 4038 -960 4150 326
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9692 354 9720 327655
rect 17960 177336 18012 177342
rect 17960 177278 18012 177284
rect 13544 13116 13596 13122
rect 13544 13058 13596 13064
rect 11888 10328 11940 10334
rect 11888 10270 11940 10276
rect 11152 7744 11204 7750
rect 11152 7686 11204 7692
rect 11164 480 11192 7686
rect 9926 354 10038 480
rect 9692 326 10038 354
rect 9926 -960 10038 326
rect 11122 -960 11234 480
rect 11900 354 11928 10270
rect 13556 480 13584 13058
rect 17038 8936 17094 8945
rect 17038 8871 17094 8880
rect 14740 4888 14792 4894
rect 14740 4830 14792 4836
rect 14752 480 14780 4830
rect 15936 3460 15988 3466
rect 15936 3402 15988 3408
rect 15948 480 15976 3402
rect 17052 480 17080 8871
rect 12318 354 12430 480
rect 11900 326 12430 354
rect 12318 -960 12430 326
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 17972 354 18000 177278
rect 24872 16574 24900 333231
rect 24872 16546 25360 16574
rect 22558 13152 22614 13161
rect 22558 13087 22614 13096
rect 20168 10532 20220 10538
rect 20168 10474 20220 10480
rect 19432 6180 19484 6186
rect 19432 6122 19484 6128
rect 19444 480 19472 6122
rect 18206 354 18318 480
rect 17972 326 18318 354
rect 18206 -960 18318 326
rect 19402 -960 19514 480
rect 20180 354 20208 10474
rect 21822 9072 21878 9081
rect 21822 9007 21878 9016
rect 21836 480 21864 9007
rect 20598 354 20710 480
rect 20180 326 20710 354
rect 20598 -960 20710 326
rect 21794 -960 21906 480
rect 22572 354 22600 13087
rect 24214 3360 24270 3369
rect 24214 3295 24270 3304
rect 24228 480 24256 3295
rect 25332 480 25360 16546
rect 22990 354 23102 480
rect 22572 326 23102 354
rect 22990 -960 23102 326
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26252 354 26280 337214
rect 52460 334552 52512 334558
rect 52460 334494 52512 334500
rect 41420 333260 41472 333266
rect 41420 333202 41472 333208
rect 34520 331900 34572 331906
rect 34520 331842 34572 331848
rect 30380 153876 30432 153882
rect 30380 153818 30432 153824
rect 27618 79384 27674 79393
rect 27618 79319 27674 79328
rect 27632 16574 27660 79319
rect 30392 16574 30420 153818
rect 27632 16546 27752 16574
rect 30392 16546 30880 16574
rect 27724 480 27752 16546
rect 28908 7812 28960 7818
rect 28908 7754 28960 7760
rect 28920 480 28948 7754
rect 30104 3528 30156 3534
rect 30104 3470 30156 3476
rect 30116 480 30144 3470
rect 26486 354 26598 480
rect 26252 326 26598 354
rect 26486 -960 26598 326
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 30852 354 30880 16546
rect 33600 11756 33652 11762
rect 33600 11698 33652 11704
rect 32402 9208 32458 9217
rect 32402 9143 32458 9152
rect 32416 480 32444 9143
rect 33612 480 33640 11698
rect 31270 354 31382 480
rect 30852 326 31382 354
rect 31270 -960 31382 326
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34532 354 34560 331842
rect 37280 329112 37332 329118
rect 37280 329054 37332 329060
rect 37292 16574 37320 329054
rect 41432 16574 41460 333202
rect 45558 331800 45614 331809
rect 45558 331735 45614 331744
rect 44180 160744 44232 160750
rect 44180 160686 44232 160692
rect 37292 16546 38424 16574
rect 41432 16546 41920 16574
rect 36728 10396 36780 10402
rect 36728 10338 36780 10344
rect 35992 8968 36044 8974
rect 35992 8910 36044 8916
rect 36004 480 36032 8910
rect 34766 354 34878 480
rect 34532 326 34878 354
rect 34766 -960 34878 326
rect 35962 -960 36074 480
rect 36740 354 36768 10338
rect 38396 480 38424 16546
rect 40222 13288 40278 13297
rect 40222 13223 40278 13232
rect 39578 9344 39634 9353
rect 39578 9279 39634 9288
rect 39592 480 39620 9279
rect 37158 354 37270 480
rect 36740 326 37270 354
rect 37158 -960 37270 326
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40236 354 40264 13223
rect 41892 480 41920 16546
rect 42800 10600 42852 10606
rect 42800 10542 42852 10548
rect 40654 354 40766 480
rect 40236 326 40766 354
rect 40654 -960 40766 326
rect 41850 -960 41962 480
rect 42812 354 42840 10542
rect 44192 3398 44220 160686
rect 45572 16574 45600 331735
rect 46940 327752 46992 327758
rect 46940 327694 46992 327700
rect 46952 16574 46980 327694
rect 49700 178764 49752 178770
rect 49700 178706 49752 178712
rect 48320 177404 48372 177410
rect 48320 177346 48372 177352
rect 48332 16574 48360 177346
rect 49712 16574 49740 178706
rect 45572 16546 46704 16574
rect 46952 16546 47440 16574
rect 48332 16546 48544 16574
rect 49712 16546 50200 16574
rect 44270 13424 44326 13433
rect 44270 13359 44326 13368
rect 44180 3392 44232 3398
rect 44180 3334 44232 3340
rect 44284 480 44312 13359
rect 45100 3392 45152 3398
rect 45100 3334 45152 3340
rect 43046 354 43158 480
rect 42812 326 43158 354
rect 43046 -960 43158 326
rect 44242 -960 44354 480
rect 45112 354 45140 3334
rect 46676 480 46704 16546
rect 45438 354 45550 480
rect 45112 326 45550 354
rect 45438 -960 45550 326
rect 46634 -960 46746 480
rect 47412 354 47440 16546
rect 47830 354 47942 480
rect 47412 326 47942 354
rect 48516 354 48544 16546
rect 50172 480 50200 16546
rect 51356 7608 51408 7614
rect 51356 7550 51408 7556
rect 51368 480 51396 7550
rect 52472 6914 52500 334494
rect 74540 331968 74592 331974
rect 74540 331910 74592 331916
rect 60740 330540 60792 330546
rect 60740 330482 60792 330488
rect 52552 329180 52604 329186
rect 52552 329122 52604 329128
rect 52564 16574 52592 329122
rect 57978 329080 58034 329089
rect 57978 329015 58034 329024
rect 55220 177472 55272 177478
rect 55220 177414 55272 177420
rect 55232 16574 55260 177414
rect 57992 16574 58020 329015
rect 52564 16546 53328 16574
rect 55232 16546 56088 16574
rect 57992 16546 58480 16574
rect 52472 6886 52592 6914
rect 52564 480 52592 6886
rect 48934 354 49046 480
rect 48516 326 49046 354
rect 47830 -960 47942 326
rect 48934 -960 49046 326
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53300 354 53328 16546
rect 54942 9480 54998 9489
rect 54942 9415 54998 9424
rect 54956 480 54984 9415
rect 56060 480 56088 16546
rect 57244 4956 57296 4962
rect 57244 4898 57296 4904
rect 57256 480 57284 4898
rect 58452 480 58480 16546
rect 59358 13560 59414 13569
rect 59358 13495 59414 13504
rect 53718 354 53830 480
rect 53300 326 53830 354
rect 53718 -960 53830 326
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59372 354 59400 13495
rect 60752 6914 60780 330482
rect 60830 329216 60886 329225
rect 60830 329151 60886 329160
rect 60844 16574 60872 329151
rect 67640 178832 67692 178838
rect 67640 178774 67692 178780
rect 66260 177540 66312 177546
rect 66260 177482 66312 177488
rect 62118 177304 62174 177313
rect 62118 177239 62174 177248
rect 62132 16574 62160 177239
rect 66272 16574 66300 177482
rect 60844 16546 61608 16574
rect 62132 16546 63264 16574
rect 66272 16546 66760 16574
rect 60752 6886 60872 6914
rect 60844 480 60872 6886
rect 59606 354 59718 480
rect 59372 326 59718 354
rect 59606 -960 59718 326
rect 60802 -960 60914 480
rect 61580 354 61608 16546
rect 63236 480 63264 16546
rect 64328 5024 64380 5030
rect 64328 4966 64380 4972
rect 64340 480 64368 4966
rect 65524 3664 65576 3670
rect 65524 3606 65576 3612
rect 65536 480 65564 3606
rect 66732 480 66760 16546
rect 61998 354 62110 480
rect 61580 326 62110 354
rect 61998 -960 62110 326
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67652 354 67680 178774
rect 74552 16574 74580 331910
rect 80058 80744 80114 80753
rect 80058 80679 80114 80688
rect 80072 16574 80100 80679
rect 81452 16574 81480 337282
rect 84200 333328 84252 333334
rect 84200 333270 84252 333276
rect 74552 16546 75040 16574
rect 80072 16546 80928 16574
rect 81452 16546 81664 16574
rect 73344 11824 73396 11830
rect 73344 11766 73396 11772
rect 69112 10464 69164 10470
rect 69112 10406 69164 10412
rect 69124 480 69152 10406
rect 72608 6248 72660 6254
rect 71502 6216 71558 6225
rect 72608 6190 72660 6196
rect 71502 6151 71558 6160
rect 70308 3800 70360 3806
rect 70308 3742 70360 3748
rect 70320 480 70348 3742
rect 71516 480 71544 6151
rect 72620 480 72648 6190
rect 67886 354 67998 480
rect 67652 326 67998 354
rect 67886 -960 67998 326
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73356 354 73384 11766
rect 75012 480 75040 16546
rect 77390 14512 77446 14521
rect 77390 14447 77446 14456
rect 75918 10296 75974 10305
rect 75918 10231 75974 10240
rect 73774 354 73886 480
rect 73356 326 73886 354
rect 73774 -960 73886 326
rect 74970 -960 75082 480
rect 75932 354 75960 10231
rect 77404 480 77432 14447
rect 79230 10432 79286 10441
rect 79230 10367 79286 10376
rect 78588 6316 78640 6322
rect 78588 6258 78640 6264
rect 78600 480 78628 6258
rect 76166 354 76278 480
rect 75932 326 76278 354
rect 76166 -960 76278 326
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79244 354 79272 10367
rect 80900 480 80928 16546
rect 79662 354 79774 480
rect 79244 326 79774 354
rect 79662 -960 79774 326
rect 80858 -960 80970 480
rect 81636 354 81664 16546
rect 83280 7676 83332 7682
rect 83280 7618 83332 7624
rect 83292 480 83320 7618
rect 82054 354 82166 480
rect 81636 326 82166 354
rect 82054 -960 82166 326
rect 83250 -960 83362 480
rect 84212 354 84240 333270
rect 90376 85542 90404 382599
rect 94504 382560 94556 382566
rect 94504 382502 94556 382508
rect 91744 382492 91796 382498
rect 91744 382434 91796 382440
rect 90456 381132 90508 381138
rect 90456 381074 90508 381080
rect 90468 241466 90496 381074
rect 91100 333396 91152 333402
rect 91100 333338 91152 333344
rect 90456 241460 90508 241466
rect 90456 241402 90508 241408
rect 90456 126268 90508 126274
rect 90456 126210 90508 126216
rect 90364 85536 90416 85542
rect 90364 85478 90416 85484
rect 86960 82136 87012 82142
rect 86960 82078 87012 82084
rect 86972 16574 87000 82078
rect 90468 33114 90496 126210
rect 90456 33108 90508 33114
rect 90456 33050 90508 33056
rect 91112 16574 91140 333338
rect 91756 255270 91784 382434
rect 93858 333432 93914 333441
rect 93858 333367 93914 333376
rect 91744 255264 91796 255270
rect 91744 255206 91796 255212
rect 92480 89004 92532 89010
rect 92480 88946 92532 88952
rect 86972 16546 87552 16574
rect 91112 16546 91600 16574
rect 85672 7880 85724 7886
rect 85672 7822 85724 7828
rect 85684 480 85712 7822
rect 86868 3732 86920 3738
rect 86868 3674 86920 3680
rect 86880 480 86908 3674
rect 84446 354 84558 480
rect 84212 326 84558 354
rect 84446 -960 84558 326
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87524 354 87552 16546
rect 89904 11960 89956 11966
rect 89904 11902 89956 11908
rect 89166 6352 89222 6361
rect 89166 6287 89222 6296
rect 89180 480 89208 6287
rect 87942 354 88054 480
rect 87524 326 88054 354
rect 87942 -960 88054 326
rect 89138 -960 89250 480
rect 89916 354 89944 11902
rect 91572 480 91600 16546
rect 90334 354 90446 480
rect 89916 326 90446 354
rect 90334 -960 90446 326
rect 91530 -960 91642 480
rect 92492 354 92520 88946
rect 93872 16574 93900 333367
rect 94516 150414 94544 382502
rect 139400 337408 139452 337414
rect 139400 337350 139452 337356
rect 128360 336116 128412 336122
rect 128360 336058 128412 336064
rect 125600 336048 125652 336054
rect 125600 335990 125652 335996
rect 118700 333464 118752 333470
rect 118700 333406 118752 333412
rect 111798 327992 111854 328001
rect 111798 327927 111854 327936
rect 96618 327856 96674 327865
rect 96618 327791 96674 327800
rect 94504 150408 94556 150414
rect 94504 150350 94556 150356
rect 96632 16574 96660 327791
rect 109040 179036 109092 179042
rect 109040 178978 109092 178984
rect 104900 178968 104952 178974
rect 104900 178910 104952 178916
rect 98000 178900 98052 178906
rect 98000 178842 98052 178848
rect 98012 16574 98040 178842
rect 99380 89072 99432 89078
rect 99380 89014 99432 89020
rect 99392 16574 99420 89014
rect 104912 16574 104940 178910
rect 93872 16546 93992 16574
rect 96632 16546 97488 16574
rect 98012 16546 98224 16574
rect 99392 16546 99880 16574
rect 104912 16546 105768 16574
rect 93964 480 93992 16546
rect 96250 7576 96306 7585
rect 96250 7511 96306 7520
rect 95146 4992 95202 5001
rect 95146 4927 95202 4936
rect 95160 480 95188 4927
rect 96264 480 96292 7511
rect 97460 480 97488 16546
rect 92726 354 92838 480
rect 92492 326 92838 354
rect 92726 -960 92838 326
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98196 354 98224 16546
rect 99852 480 99880 16546
rect 102232 14476 102284 14482
rect 102232 14418 102284 14424
rect 100760 12028 100812 12034
rect 100760 11970 100812 11976
rect 98614 354 98726 480
rect 98196 326 98726 354
rect 98614 -960 98726 326
rect 99810 -960 99922 480
rect 100772 354 100800 11970
rect 102244 480 102272 14418
rect 104072 12096 104124 12102
rect 104072 12038 104124 12044
rect 103336 7948 103388 7954
rect 103336 7890 103388 7896
rect 103348 480 103376 7890
rect 101006 354 101118 480
rect 100772 326 101118 354
rect 101006 -960 101118 326
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104084 354 104112 12038
rect 105740 480 105768 16546
rect 108120 12164 108172 12170
rect 108120 12106 108172 12112
rect 106924 9036 106976 9042
rect 106924 8978 106976 8984
rect 106936 480 106964 8978
rect 108132 480 108160 12106
rect 104502 354 104614 480
rect 104084 326 104614 354
rect 104502 -960 104614 326
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109052 354 109080 178978
rect 111812 16574 111840 327927
rect 115940 179104 115992 179110
rect 115940 179046 115992 179052
rect 114558 44840 114614 44849
rect 114558 44775 114614 44784
rect 114572 16574 114600 44775
rect 115952 16574 115980 179046
rect 118712 16574 118740 333406
rect 122840 332036 122892 332042
rect 122840 331978 122892 331984
rect 122852 16574 122880 331978
rect 111812 16546 112392 16574
rect 114572 16546 114784 16574
rect 115952 16546 116440 16574
rect 118712 16546 118832 16574
rect 122852 16546 123064 16574
rect 110512 14544 110564 14550
rect 110512 14486 110564 14492
rect 110524 480 110552 14486
rect 111614 13696 111670 13705
rect 111614 13631 111670 13640
rect 111628 480 111656 13631
rect 109286 354 109398 480
rect 109052 326 109398 354
rect 109286 -960 109398 326
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112364 354 112392 16546
rect 114008 10668 114060 10674
rect 114008 10610 114060 10616
rect 114020 480 114048 10610
rect 112782 354 112894 480
rect 112364 326 112894 354
rect 112782 -960 112894 326
rect 113978 -960 114090 480
rect 114756 354 114784 16546
rect 116412 480 116440 16546
rect 117320 12232 117372 12238
rect 117320 12174 117372 12180
rect 115174 354 115286 480
rect 114756 326 115286 354
rect 115174 -960 115286 326
rect 116370 -960 116482 480
rect 117332 354 117360 12174
rect 118804 480 118832 16546
rect 120632 14612 120684 14618
rect 120632 14554 120684 14560
rect 119894 6488 119950 6497
rect 119894 6423 119950 6432
rect 119908 480 119936 6423
rect 117566 354 117678 480
rect 117332 326 117678 354
rect 117566 -960 117678 326
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 120644 354 120672 14554
rect 122288 13184 122340 13190
rect 122288 13126 122340 13132
rect 122300 480 122328 13126
rect 121062 354 121174 480
rect 120644 326 121174 354
rect 121062 -960 121174 326
rect 122258 -960 122370 480
rect 123036 354 123064 16546
rect 124680 13252 124732 13258
rect 124680 13194 124732 13200
rect 124692 480 124720 13194
rect 123454 354 123566 480
rect 123036 326 123566 354
rect 123454 -960 123566 326
rect 124650 -960 124762 480
rect 125612 354 125640 335990
rect 126980 329248 127032 329254
rect 126980 329190 127032 329196
rect 126992 480 127020 329190
rect 128372 16574 128400 336058
rect 136640 334756 136692 334762
rect 136640 334698 136692 334704
rect 133880 334688 133932 334694
rect 133880 334630 133932 334636
rect 132498 330440 132554 330449
rect 132498 330375 132554 330384
rect 129738 326496 129794 326505
rect 129738 326431 129794 326440
rect 129752 16574 129780 326431
rect 132512 16574 132540 330375
rect 128372 16546 128952 16574
rect 129752 16546 130608 16574
rect 132512 16546 133000 16574
rect 127624 12300 127676 12306
rect 127624 12242 127676 12248
rect 127636 3806 127664 12242
rect 128176 3936 128228 3942
rect 128176 3878 128228 3884
rect 127624 3800 127676 3806
rect 127624 3742 127676 3748
rect 128188 480 128216 3878
rect 125846 354 125958 480
rect 125612 326 125958 354
rect 125846 -960 125958 326
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 128924 354 128952 16546
rect 130580 480 130608 16546
rect 131762 9616 131818 9625
rect 131762 9551 131818 9560
rect 131776 480 131804 9551
rect 132972 480 133000 16546
rect 129342 354 129454 480
rect 128924 326 129454 354
rect 129342 -960 129454 326
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 133892 354 133920 334630
rect 135260 333532 135312 333538
rect 135260 333474 135312 333480
rect 135272 480 135300 333474
rect 136652 16574 136680 334698
rect 139412 16574 139440 337350
rect 165620 337068 165672 337074
rect 165620 337010 165672 337016
rect 161480 337000 161532 337006
rect 161480 336942 161532 336948
rect 160100 336184 160152 336190
rect 160100 336126 160152 336132
rect 151820 334824 151872 334830
rect 151820 334766 151872 334772
rect 147678 334656 147734 334665
rect 147678 334591 147734 334600
rect 146298 330576 146354 330585
rect 146298 330511 146354 330520
rect 144920 177608 144972 177614
rect 144920 177550 144972 177556
rect 142160 21412 142212 21418
rect 142160 21354 142212 21360
rect 136652 16546 137232 16574
rect 139412 16546 139624 16574
rect 136454 3496 136510 3505
rect 136454 3431 136510 3440
rect 136468 480 136496 3431
rect 134126 354 134238 480
rect 133892 326 134238 354
rect 134126 -960 134238 326
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137204 354 137232 16546
rect 138848 9104 138900 9110
rect 138848 9046 138900 9052
rect 138860 480 138888 9046
rect 137622 354 137734 480
rect 137204 326 137734 354
rect 137622 -960 137734 326
rect 138818 -960 138930 480
rect 139596 354 139624 16546
rect 141240 3868 141292 3874
rect 141240 3810 141292 3816
rect 141252 480 141280 3810
rect 140014 354 140126 480
rect 139596 326 140126 354
rect 140014 -960 140126 326
rect 141210 -960 141322 480
rect 142172 354 142200 21354
rect 144932 16574 144960 177550
rect 146312 16574 146340 330511
rect 147692 16574 147720 334591
rect 149060 333872 149112 333878
rect 149060 333814 149112 333820
rect 149072 16574 149100 333814
rect 150438 328128 150494 328137
rect 150438 328063 150494 328072
rect 150452 16574 150480 328063
rect 144932 16546 145512 16574
rect 146312 16546 147168 16574
rect 147692 16546 147904 16574
rect 149072 16546 149560 16574
rect 150452 16546 150664 16574
rect 143540 8016 143592 8022
rect 143540 7958 143592 7964
rect 143552 480 143580 7958
rect 144734 6624 144790 6633
rect 144734 6559 144790 6568
rect 144748 480 144776 6559
rect 142406 354 142518 480
rect 142172 326 142518 354
rect 142406 -960 142518 326
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145484 354 145512 16546
rect 147140 480 147168 16546
rect 145902 354 146014 480
rect 145484 326 146014 354
rect 145902 -960 146014 326
rect 147098 -960 147210 480
rect 147876 354 147904 16546
rect 149532 480 149560 16546
rect 150636 480 150664 16546
rect 151832 480 151860 334766
rect 155960 333668 156012 333674
rect 155960 333610 156012 333616
rect 153200 329316 153252 329322
rect 153200 329258 153252 329264
rect 151912 177676 151964 177682
rect 151912 177618 151964 177624
rect 151924 16574 151952 177618
rect 153212 16574 153240 329258
rect 154580 191140 154632 191146
rect 154580 191082 154632 191088
rect 154592 16574 154620 191082
rect 155972 16574 156000 333610
rect 158720 177744 158772 177750
rect 158720 177686 158772 177692
rect 158732 16574 158760 177686
rect 151924 16546 153056 16574
rect 153212 16546 153792 16574
rect 154592 16546 155448 16574
rect 155972 16546 156184 16574
rect 158732 16546 158944 16574
rect 153028 480 153056 16546
rect 148294 354 148406 480
rect 147876 326 148406 354
rect 148294 -960 148406 326
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 153764 354 153792 16546
rect 155420 480 155448 16546
rect 154182 354 154294 480
rect 153764 326 154294 354
rect 154182 -960 154294 326
rect 155378 -960 155490 480
rect 156156 354 156184 16546
rect 157798 5128 157854 5137
rect 157798 5063 157854 5072
rect 157812 480 157840 5063
rect 158916 480 158944 16546
rect 160112 11694 160140 336126
rect 160192 179172 160244 179178
rect 160192 179114 160244 179120
rect 160100 11688 160152 11694
rect 160100 11630 160152 11636
rect 160204 6914 160232 179114
rect 161492 16574 161520 336942
rect 164238 336016 164294 336025
rect 164238 335951 164294 335960
rect 162860 177812 162912 177818
rect 162860 177754 162912 177760
rect 162872 16574 162900 177754
rect 164252 16574 164280 335951
rect 165632 16574 165660 337010
rect 173900 334892 173952 334898
rect 173900 334834 173952 334840
rect 168380 332104 168432 332110
rect 168380 332046 168432 332052
rect 161492 16546 162072 16574
rect 162872 16546 163728 16574
rect 164252 16546 164464 16574
rect 165632 16546 166120 16574
rect 161296 11688 161348 11694
rect 161296 11630 161348 11636
rect 160112 6886 160232 6914
rect 160112 480 160140 6886
rect 161308 480 161336 11630
rect 156574 354 156686 480
rect 156156 326 156686 354
rect 156574 -960 156686 326
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162044 354 162072 16546
rect 163700 480 163728 16546
rect 162462 354 162574 480
rect 162044 326 162574 354
rect 162462 -960 162574 326
rect 163658 -960 163770 480
rect 164436 354 164464 16546
rect 166092 480 166120 16546
rect 167182 7712 167238 7721
rect 167182 7647 167238 7656
rect 167196 480 167224 7647
rect 168392 480 168420 332046
rect 171140 327820 171192 327826
rect 171140 327762 171192 327768
rect 171152 16574 171180 327762
rect 171152 16546 172008 16574
rect 170772 8084 170824 8090
rect 170772 8026 170824 8032
rect 169574 6760 169630 6769
rect 169574 6695 169630 6704
rect 169588 480 169616 6695
rect 170784 480 170812 8026
rect 171980 480 172008 16546
rect 173164 6384 173216 6390
rect 173164 6326 173216 6332
rect 173176 480 173204 6326
rect 164854 354 164966 480
rect 164436 326 164966 354
rect 164854 -960 164966 326
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 173912 354 173940 334834
rect 174556 20670 174584 384610
rect 231124 384260 231176 384266
rect 231124 384202 231176 384208
rect 174636 382628 174688 382634
rect 174636 382570 174688 382576
rect 174648 372570 174676 382570
rect 174636 372564 174688 372570
rect 174636 372506 174688 372512
rect 227720 337204 227772 337210
rect 227720 337146 227772 337152
rect 218060 337136 218112 337142
rect 218060 337078 218112 337084
rect 196624 336456 196676 336462
rect 182822 336424 182878 336433
rect 196624 336398 196676 336404
rect 182822 336359 182878 336368
rect 178866 336288 178922 336297
rect 178866 336223 178922 336232
rect 182180 336252 182232 336258
rect 178682 336152 178738 336161
rect 178682 336087 178738 336096
rect 176660 177880 176712 177886
rect 176660 177822 176712 177828
rect 174544 20664 174596 20670
rect 174544 20606 174596 20612
rect 175924 5092 175976 5098
rect 175924 5034 175976 5040
rect 175464 3800 175516 3806
rect 175464 3742 175516 3748
rect 175476 480 175504 3742
rect 175936 3602 175964 5034
rect 175924 3596 175976 3602
rect 175924 3538 175976 3544
rect 176672 480 176700 177822
rect 176752 159384 176804 159390
rect 176752 159326 176804 159332
rect 176764 16574 176792 159326
rect 176764 16546 177896 16574
rect 177868 480 177896 16546
rect 178696 7750 178724 336087
rect 178880 11898 178908 336223
rect 182180 336194 182232 336200
rect 180800 327888 180852 327894
rect 180800 327830 180852 327836
rect 180812 16574 180840 327830
rect 180812 16546 181024 16574
rect 178868 11892 178920 11898
rect 178868 11834 178920 11840
rect 178684 7744 178736 7750
rect 178684 7686 178736 7692
rect 180248 7744 180300 7750
rect 180248 7686 180300 7692
rect 179052 3596 179104 3602
rect 179052 3538 179104 3544
rect 179064 480 179092 3538
rect 180260 480 180288 7686
rect 174238 354 174350 480
rect 173912 326 174350 354
rect 174238 -960 174350 326
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 180996 354 181024 16546
rect 181444 10736 181496 10742
rect 181444 10678 181496 10684
rect 181456 3738 181484 10678
rect 181444 3732 181496 3738
rect 181444 3674 181496 3680
rect 181414 354 181526 480
rect 180996 326 181526 354
rect 182192 354 182220 336194
rect 182836 10538 182864 336359
rect 188344 336320 188396 336326
rect 188344 336262 188396 336268
rect 184940 330676 184992 330682
rect 184940 330618 184992 330624
rect 183558 326632 183614 326641
rect 183558 326567 183614 326576
rect 183572 16574 183600 326567
rect 183572 16546 183784 16574
rect 182824 10532 182876 10538
rect 182824 10474 182876 10480
rect 182914 6896 182970 6905
rect 182914 6831 182970 6840
rect 182928 3942 182956 6831
rect 182916 3936 182968 3942
rect 182916 3878 182968 3884
rect 183756 480 183784 16546
rect 184952 11694 184980 330618
rect 187700 158024 187752 158030
rect 187700 157966 187752 157972
rect 186318 155408 186374 155417
rect 186318 155343 186374 155352
rect 185030 155272 185086 155281
rect 185030 155207 185086 155216
rect 184940 11688 184992 11694
rect 184940 11630 184992 11636
rect 185044 6914 185072 155207
rect 186332 16574 186360 155343
rect 186332 16546 186912 16574
rect 186136 11688 186188 11694
rect 186136 11630 186188 11636
rect 184952 6886 185072 6914
rect 184952 480 184980 6886
rect 186148 480 186176 11630
rect 182518 354 182630 480
rect 182192 326 182630 354
rect 181414 -960 181526 326
rect 182518 -960 182630 326
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 186884 354 186912 16546
rect 187712 6914 187740 157966
rect 188356 7818 188384 336262
rect 193220 330744 193272 330750
rect 193220 330686 193272 330692
rect 189080 330608 189132 330614
rect 189080 330550 189132 330556
rect 189092 16574 189120 330550
rect 191840 320884 191892 320890
rect 191840 320826 191892 320832
rect 190460 155236 190512 155242
rect 190460 155178 190512 155184
rect 189092 16546 189304 16574
rect 188344 7812 188396 7818
rect 188344 7754 188396 7760
rect 187712 6886 188568 6914
rect 188540 480 188568 6886
rect 187302 354 187414 480
rect 186884 326 187414 354
rect 187302 -960 187414 326
rect 188498 -960 188610 480
rect 189276 354 189304 16546
rect 189694 354 189806 480
rect 189276 326 189806 354
rect 190472 354 190500 155178
rect 191852 16574 191880 320826
rect 191852 16546 192064 16574
rect 192036 480 192064 16546
rect 193232 480 193260 330686
rect 194600 155372 194652 155378
rect 194600 155314 194652 155320
rect 193312 155304 193364 155310
rect 193312 155246 193364 155252
rect 193324 16574 193352 155246
rect 194612 16574 194640 155314
rect 193324 16546 194456 16574
rect 194612 16546 195192 16574
rect 194428 480 194456 16546
rect 190798 354 190910 480
rect 190472 326 190910 354
rect 189694 -960 189806 326
rect 190798 -960 190910 326
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195164 354 195192 16546
rect 196072 9580 196124 9586
rect 196072 9522 196124 9528
rect 196084 3670 196112 9522
rect 196636 8974 196664 336398
rect 200764 336388 200816 336394
rect 200764 336330 200816 336336
rect 197360 155440 197412 155446
rect 197360 155382 197412 155388
rect 197372 16574 197400 155382
rect 197372 16546 197952 16574
rect 196624 8968 196676 8974
rect 196624 8910 196676 8916
rect 197360 5160 197412 5166
rect 197360 5102 197412 5108
rect 197372 3874 197400 5102
rect 197360 3868 197412 3874
rect 197360 3810 197412 3816
rect 196808 3732 196860 3738
rect 196808 3674 196860 3680
rect 196072 3664 196124 3670
rect 196072 3606 196124 3612
rect 196820 480 196848 3674
rect 197924 480 197952 16546
rect 200776 10606 200804 336330
rect 211160 334960 211212 334966
rect 211160 334902 211212 334908
rect 207020 330812 207072 330818
rect 207020 330754 207072 330760
rect 204260 158092 204312 158098
rect 204260 158034 204312 158040
rect 201498 156632 201554 156641
rect 201498 156567 201554 156576
rect 201512 11694 201540 156567
rect 201590 155544 201646 155553
rect 201590 155479 201646 155488
rect 201500 11688 201552 11694
rect 201500 11630 201552 11636
rect 200764 10600 200816 10606
rect 200764 10542 200816 10548
rect 199108 7812 199160 7818
rect 199108 7754 199160 7760
rect 199120 480 199148 7754
rect 201604 6914 201632 155479
rect 204272 16574 204300 158034
rect 205640 156664 205692 156670
rect 205640 156606 205692 156612
rect 205652 16574 205680 156606
rect 204272 16546 205128 16574
rect 205652 16546 206232 16574
rect 202696 11688 202748 11694
rect 202696 11630 202748 11636
rect 201512 6886 201632 6914
rect 200304 3664 200356 3670
rect 200304 3606 200356 3612
rect 200316 480 200344 3606
rect 201512 480 201540 6886
rect 202708 480 202736 11630
rect 203892 3868 203944 3874
rect 203892 3810 203944 3816
rect 203904 480 203932 3810
rect 205100 480 205128 16546
rect 206204 480 206232 16546
rect 195582 354 195694 480
rect 195164 326 195694 354
rect 195582 -960 195694 326
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207032 354 207060 330754
rect 209780 326392 209832 326398
rect 209780 326334 209832 326340
rect 208400 158160 208452 158166
rect 208400 158102 208452 158108
rect 208412 16574 208440 158102
rect 208412 16546 208624 16574
rect 208596 480 208624 16546
rect 209792 480 209820 326334
rect 209870 155680 209926 155689
rect 209870 155615 209926 155624
rect 209884 16574 209912 155615
rect 211172 16574 211200 334902
rect 216680 333736 216732 333742
rect 216680 333678 216732 333684
rect 215298 160712 215354 160721
rect 215298 160647 215354 160656
rect 212540 159452 212592 159458
rect 212540 159394 212592 159400
rect 212552 16574 212580 159394
rect 213920 156732 213972 156738
rect 213920 156674 213972 156680
rect 213932 16574 213960 156674
rect 209884 16546 211016 16574
rect 211172 16546 211752 16574
rect 212552 16546 213408 16574
rect 213932 16546 214512 16574
rect 210988 480 211016 16546
rect 207358 354 207470 480
rect 207032 326 207470 354
rect 207358 -960 207470 326
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 211724 354 211752 16546
rect 213380 480 213408 16546
rect 214484 480 214512 16546
rect 212142 354 212254 480
rect 211724 326 212254 354
rect 212142 -960 212254 326
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215312 354 215340 160647
rect 216692 16574 216720 333678
rect 216692 16546 216904 16574
rect 216876 480 216904 16546
rect 218072 480 218100 337078
rect 224960 336524 225012 336530
rect 224960 336466 225012 336472
rect 220820 329384 220872 329390
rect 220820 329326 220872 329332
rect 219440 158228 219492 158234
rect 219440 158170 219492 158176
rect 218150 157992 218206 158001
rect 218150 157927 218206 157936
rect 218164 16574 218192 157927
rect 219452 16574 219480 158170
rect 220832 16574 220860 329326
rect 223580 159588 223632 159594
rect 223580 159530 223632 159536
rect 222200 159520 222252 159526
rect 222200 159462 222252 159468
rect 222212 16574 222240 159462
rect 218164 16546 219296 16574
rect 219452 16546 220032 16574
rect 220832 16546 221136 16574
rect 222212 16546 222792 16574
rect 219268 480 219296 16546
rect 215638 354 215750 480
rect 215312 326 215750 354
rect 215638 -960 215750 326
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220004 354 220032 16546
rect 220422 354 220534 480
rect 220004 326 220534 354
rect 221108 354 221136 16546
rect 221464 10532 221516 10538
rect 221464 10474 221516 10480
rect 221476 3534 221504 10474
rect 221464 3528 221516 3534
rect 221464 3470 221516 3476
rect 222764 480 222792 16546
rect 221526 354 221638 480
rect 221108 326 221638 354
rect 220422 -960 220534 326
rect 221526 -960 221638 326
rect 222722 -960 222834 480
rect 223592 354 223620 159530
rect 224972 16574 225000 336466
rect 226340 332308 226392 332314
rect 226340 332250 226392 332256
rect 224972 16546 225184 16574
rect 225156 480 225184 16546
rect 226352 3534 226380 332250
rect 227732 16574 227760 337146
rect 229100 335028 229152 335034
rect 229100 334970 229152 334976
rect 229112 16574 229140 334970
rect 230480 159656 230532 159662
rect 230480 159598 230532 159604
rect 230492 16574 230520 159598
rect 231136 59362 231164 384202
rect 233976 383988 234028 383994
rect 233976 383930 234028 383936
rect 233792 382424 233844 382430
rect 233792 382366 233844 382372
rect 232504 382288 232556 382294
rect 232504 382230 232556 382236
rect 232516 267034 232544 382230
rect 233240 335096 233292 335102
rect 233240 335038 233292 335044
rect 232504 267028 232556 267034
rect 232504 266970 232556 266976
rect 231860 156800 231912 156806
rect 231860 156742 231912 156748
rect 231124 59356 231176 59362
rect 231124 59298 231176 59304
rect 227732 16546 228312 16574
rect 229112 16546 229416 16574
rect 230492 16546 231072 16574
rect 226340 3528 226392 3534
rect 226340 3470 226392 3476
rect 227536 3528 227588 3534
rect 227536 3470 227588 3476
rect 227628 3528 227680 3534
rect 227628 3470 227680 3476
rect 226340 2848 226392 2854
rect 226340 2790 226392 2796
rect 226352 480 226380 2790
rect 227548 480 227576 3470
rect 227640 2854 227668 3470
rect 227628 2848 227680 2854
rect 227628 2790 227680 2796
rect 223918 354 224030 480
rect 223592 326 224030 354
rect 223918 -960 224030 326
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228284 354 228312 16546
rect 228702 354 228814 480
rect 228284 326 228814 354
rect 229388 354 229416 16546
rect 231044 480 231072 16546
rect 229806 354 229918 480
rect 229388 326 229918 354
rect 228702 -960 228814 326
rect 229806 -960 229918 326
rect 231002 -960 231114 480
rect 231872 354 231900 156742
rect 232516 131102 232544 266970
rect 232504 131096 232556 131102
rect 232504 131038 232556 131044
rect 233252 16574 233280 335038
rect 233804 306338 233832 382366
rect 233884 332240 233936 332246
rect 233884 332182 233936 332188
rect 233792 306332 233844 306338
rect 233792 306274 233844 306280
rect 233252 16546 233464 16574
rect 233436 480 233464 16546
rect 233896 3602 233924 332182
rect 233988 153202 234016 383930
rect 234080 158409 234108 389422
rect 234160 382832 234212 382838
rect 234160 382774 234212 382780
rect 234066 158400 234122 158409
rect 234066 158335 234122 158344
rect 233976 153196 234028 153202
rect 233976 153138 234028 153144
rect 234172 144906 234200 382774
rect 234252 382764 234304 382770
rect 234252 382706 234304 382712
rect 234160 144900 234212 144906
rect 234160 144842 234212 144848
rect 234264 135250 234292 382706
rect 234436 381268 234488 381274
rect 234436 381210 234488 381216
rect 234342 380488 234398 380497
rect 234342 380423 234398 380432
rect 234252 135244 234304 135250
rect 234252 135186 234304 135192
rect 234356 113150 234384 380423
rect 234344 113144 234396 113150
rect 234344 113086 234396 113092
rect 234448 97578 234476 381210
rect 234540 104854 234568 409838
rect 234632 387462 234660 703582
rect 235000 703474 235028 703582
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 299492 703582 299980 703610
rect 235184 703474 235212 703520
rect 235000 703446 235212 703474
rect 255596 700528 255648 700534
rect 255596 700470 255648 700476
rect 242164 700460 242216 700466
rect 242164 700402 242216 700408
rect 242176 394126 242204 700402
rect 253204 683188 253256 683194
rect 253204 683130 253256 683136
rect 251824 670744 251876 670750
rect 251824 670686 251876 670692
rect 249892 630692 249944 630698
rect 249892 630634 249944 630640
rect 249156 484424 249208 484430
rect 249156 484366 249208 484372
rect 247132 470620 247184 470626
rect 247132 470562 247184 470568
rect 245752 430636 245804 430642
rect 245752 430578 245804 430584
rect 242164 394120 242216 394126
rect 242164 394062 242216 394068
rect 234620 387456 234672 387462
rect 234620 387398 234672 387404
rect 235816 386436 235868 386442
rect 235816 386378 235868 386384
rect 235540 385892 235592 385898
rect 235540 385834 235592 385840
rect 235552 385218 235580 385834
rect 235540 385212 235592 385218
rect 235540 385154 235592 385160
rect 235724 385212 235776 385218
rect 235724 385154 235776 385160
rect 235632 384396 235684 384402
rect 235632 384338 235684 384344
rect 235448 383104 235500 383110
rect 235448 383046 235500 383052
rect 235172 382900 235224 382906
rect 235172 382842 235224 382848
rect 235184 346390 235212 382842
rect 235262 382800 235318 382809
rect 235262 382735 235318 382744
rect 235172 346384 235224 346390
rect 235172 346326 235224 346332
rect 234620 336796 234672 336802
rect 234620 336738 234672 336744
rect 234528 104848 234580 104854
rect 234528 104790 234580 104796
rect 234436 97572 234488 97578
rect 234436 97514 234488 97520
rect 234632 11694 234660 336738
rect 234712 330880 234764 330886
rect 234712 330822 234764 330828
rect 234620 11688 234672 11694
rect 234620 11630 234672 11636
rect 234724 6914 234752 330822
rect 234804 164212 234856 164218
rect 234804 164154 234856 164160
rect 234816 163538 234844 164154
rect 234804 163532 234856 163538
rect 234804 163474 234856 163480
rect 235276 137970 235304 382735
rect 235356 382356 235408 382362
rect 235356 382298 235408 382304
rect 235368 293962 235396 382298
rect 235460 320210 235488 383046
rect 235540 381608 235592 381614
rect 235540 381550 235592 381556
rect 235448 320204 235500 320210
rect 235448 320146 235500 320152
rect 235356 293956 235408 293962
rect 235356 293898 235408 293904
rect 235552 163538 235580 381550
rect 235540 163532 235592 163538
rect 235540 163474 235592 163480
rect 235264 137964 235316 137970
rect 235264 137906 235316 137912
rect 235644 126954 235672 384338
rect 234804 126948 234856 126954
rect 234804 126890 234856 126896
rect 235632 126948 235684 126954
rect 235632 126890 235684 126896
rect 234816 126274 234844 126890
rect 234804 126268 234856 126274
rect 234804 126210 234856 126216
rect 235736 122806 235764 385154
rect 235724 122800 235776 122806
rect 235724 122742 235776 122748
rect 235828 97510 235856 386378
rect 244924 385348 244976 385354
rect 244924 385290 244976 385296
rect 244096 385076 244148 385082
rect 244096 385018 244148 385024
rect 241060 384872 241112 384878
rect 241060 384814 241112 384820
rect 236828 384804 236880 384810
rect 236828 384746 236880 384752
rect 236840 381750 236868 384746
rect 239218 384432 239274 384441
rect 239218 384367 239274 384376
rect 239232 381970 239260 384367
rect 240048 384056 240100 384062
rect 240048 383998 240100 384004
rect 239404 383784 239456 383790
rect 239404 383726 239456 383732
rect 239232 381942 239292 381970
rect 236828 381744 236880 381750
rect 236828 381686 236880 381692
rect 235908 381676 235960 381682
rect 235908 381618 235960 381624
rect 235816 97504 235868 97510
rect 235816 97446 235868 97452
rect 235920 71738 235948 381618
rect 239416 381546 239444 383726
rect 239678 381984 239734 381993
rect 239568 381942 239678 381970
rect 240060 381970 240088 383998
rect 240782 382120 240838 382129
rect 240782 382055 240838 382064
rect 240796 381970 240824 382055
rect 241072 381970 241100 384814
rect 243820 384600 243872 384606
rect 243820 384542 243872 384548
rect 242808 384532 242860 384538
rect 242808 384474 242860 384480
rect 241336 384124 241388 384130
rect 241336 384066 241388 384072
rect 241348 381970 241376 384066
rect 242162 383888 242218 383897
rect 242162 383823 242218 383832
rect 241426 382392 241482 382401
rect 241426 382327 241482 382336
rect 240060 381942 240120 381970
rect 240672 381942 240824 381970
rect 240948 381942 241100 381970
rect 241224 381942 241376 381970
rect 241440 381970 241468 382327
rect 242176 381970 242204 383823
rect 242438 383072 242494 383081
rect 242438 383007 242494 383016
rect 242452 381970 242480 383007
rect 241440 381942 241500 381970
rect 242052 381942 242204 381970
rect 242328 381942 242480 381970
rect 242820 381970 242848 384474
rect 243266 383208 243322 383217
rect 243266 383143 243322 383152
rect 243280 381970 243308 383143
rect 243832 381970 243860 384542
rect 244108 381970 244136 385018
rect 244648 383240 244700 383246
rect 244648 383182 244700 383188
rect 244660 381970 244688 383182
rect 244936 381970 244964 385290
rect 245200 383852 245252 383858
rect 245200 383794 245252 383800
rect 245212 381970 245240 383794
rect 245660 383308 245712 383314
rect 245660 383250 245712 383256
rect 245476 383172 245528 383178
rect 245476 383114 245528 383120
rect 245488 381970 245516 383114
rect 245672 382974 245700 383250
rect 245764 382974 245792 430578
rect 246028 404388 246080 404394
rect 246028 404330 246080 404336
rect 246040 402974 246068 404330
rect 246040 402946 246620 402974
rect 246396 384736 246448 384742
rect 246396 384678 246448 384684
rect 245660 382968 245712 382974
rect 245660 382910 245712 382916
rect 245752 382968 245804 382974
rect 245752 382910 245804 382916
rect 246120 382696 246172 382702
rect 246120 382638 246172 382644
rect 242820 381942 242880 381970
rect 242992 381948 243044 381954
rect 239678 381919 239734 381928
rect 243156 381942 243308 381970
rect 243708 381942 243860 381970
rect 243984 381942 244136 381970
rect 244536 381942 244688 381970
rect 244812 381942 244964 381970
rect 245088 381942 245240 381970
rect 245364 381942 245516 381970
rect 246026 381984 246082 381993
rect 246132 381970 246160 382638
rect 246302 382120 246358 382129
rect 246302 382055 246358 382064
rect 246132 381942 246192 381970
rect 246026 381919 246082 381928
rect 242992 381890 243044 381896
rect 241612 381880 241664 381886
rect 241612 381822 241664 381828
rect 239404 381540 239456 381546
rect 239404 381482 239456 381488
rect 241624 381478 241652 381822
rect 241886 381712 241942 381721
rect 241776 381670 241886 381698
rect 241886 381647 241942 381656
rect 243004 381478 243032 381890
rect 245764 381818 245916 381834
rect 245752 381812 245916 381818
rect 245804 381806 245916 381812
rect 245752 381754 245804 381760
rect 243544 381744 243596 381750
rect 243432 381692 243544 381698
rect 243432 381686 243596 381692
rect 243432 381670 243584 381686
rect 241612 381472 241664 381478
rect 239954 381440 240010 381449
rect 239844 381398 239954 381426
rect 240506 381440 240562 381449
rect 240396 381398 240506 381426
rect 239954 381375 240010 381384
rect 242992 381472 243044 381478
rect 242714 381440 242770 381449
rect 241612 381414 241664 381420
rect 242604 381398 242714 381426
rect 240506 381375 240562 381384
rect 244372 381472 244424 381478
rect 242992 381414 243044 381420
rect 244260 381420 244372 381426
rect 246040 381449 246068 381919
rect 246316 381585 246344 382055
rect 246408 381970 246436 384678
rect 246592 381970 246620 402946
rect 247144 385286 247172 470562
rect 247408 456816 247460 456822
rect 247408 456758 247460 456764
rect 247224 418192 247276 418198
rect 247224 418134 247276 418140
rect 247132 385280 247184 385286
rect 247132 385222 247184 385228
rect 246856 382968 246908 382974
rect 246856 382910 246908 382916
rect 246868 381970 246896 382910
rect 247236 381970 247264 418134
rect 247420 381970 247448 456758
rect 248512 406428 248564 406434
rect 248512 406370 248564 406376
rect 248524 392494 248552 406370
rect 248788 392624 248840 392630
rect 248788 392566 248840 392572
rect 248512 392488 248564 392494
rect 248512 392430 248564 392436
rect 248420 389836 248472 389842
rect 248420 389778 248472 389784
rect 248432 389174 248460 389778
rect 248432 389146 248552 389174
rect 248328 387320 248380 387326
rect 248328 387262 248380 387268
rect 247776 386504 247828 386510
rect 247776 386446 247828 386452
rect 247788 381970 247816 386446
rect 247960 385280 248012 385286
rect 247960 385222 248012 385228
rect 247972 381970 248000 385222
rect 248340 381970 248368 387262
rect 248524 381970 248552 389146
rect 248800 381970 248828 392566
rect 249168 386510 249196 484366
rect 249904 402974 249932 630634
rect 249904 402946 250484 402974
rect 249616 392488 249668 392494
rect 249616 392430 249668 392436
rect 249340 390108 249392 390114
rect 249340 390050 249392 390056
rect 249248 387116 249300 387122
rect 249248 387058 249300 387064
rect 249156 386504 249208 386510
rect 249156 386446 249208 386452
rect 249260 386414 249288 387058
rect 249168 386386 249288 386414
rect 248880 383920 248932 383926
rect 248880 383862 248932 383868
rect 248892 383314 248920 383862
rect 248880 383308 248932 383314
rect 248880 383250 248932 383256
rect 249064 383240 249116 383246
rect 249064 383182 249116 383188
rect 249076 382401 249104 383182
rect 249062 382392 249118 382401
rect 249062 382327 249118 382336
rect 246408 381942 246468 381970
rect 246592 381942 246744 381970
rect 246868 381942 247020 381970
rect 247236 381942 247296 381970
rect 247420 381942 247572 381970
rect 247788 381942 247848 381970
rect 247972 381942 248124 381970
rect 248236 381948 248288 381954
rect 248340 381942 248400 381970
rect 248524 381942 248676 381970
rect 248800 381942 248952 381970
rect 248236 381890 248288 381896
rect 247408 381744 247460 381750
rect 247408 381686 247460 381692
rect 247684 381744 247736 381750
rect 247684 381686 247736 381692
rect 246302 381576 246358 381585
rect 246302 381511 246358 381520
rect 247420 381478 247448 381686
rect 247696 381546 247724 381686
rect 247684 381540 247736 381546
rect 247684 381482 247736 381488
rect 248248 381478 248276 381890
rect 249168 381834 249196 386386
rect 249352 381970 249380 390050
rect 249628 381970 249656 392430
rect 250168 390176 250220 390182
rect 250168 390118 250220 390124
rect 249984 386572 250036 386578
rect 249984 386514 250036 386520
rect 249996 381970 250024 386514
rect 250180 381970 250208 390118
rect 250456 381970 250484 402946
rect 251272 392692 251324 392698
rect 251272 392634 251324 392640
rect 250996 390040 251048 390046
rect 250996 389982 251048 389988
rect 250812 386504 250864 386510
rect 250812 386446 250864 386452
rect 250824 381970 250852 386446
rect 251008 381970 251036 389982
rect 251284 385286 251312 392634
rect 251364 390584 251416 390590
rect 251364 390526 251416 390532
rect 251272 385280 251324 385286
rect 251272 385222 251324 385228
rect 251376 381970 251404 390526
rect 251640 387184 251692 387190
rect 251640 387126 251692 387132
rect 251652 381970 251680 387126
rect 251836 386510 251864 670686
rect 251916 616888 251968 616894
rect 251916 616830 251968 616836
rect 251928 386578 251956 616830
rect 252652 589960 252704 589966
rect 252652 589902 252704 589908
rect 252008 389904 252060 389910
rect 252008 389846 252060 389852
rect 251916 386572 251968 386578
rect 251916 386514 251968 386520
rect 251824 386504 251876 386510
rect 251824 386446 251876 386452
rect 252020 382242 252048 389846
rect 252468 388612 252520 388618
rect 252468 388554 252520 388560
rect 252100 385280 252152 385286
rect 252100 385222 252152 385228
rect 251974 382214 252048 382242
rect 249352 381942 249504 381970
rect 249628 381942 249780 381970
rect 249996 381942 250056 381970
rect 250180 381942 250332 381970
rect 250456 381942 250608 381970
rect 250824 381942 250884 381970
rect 251008 381942 251160 381970
rect 251376 381942 251436 381970
rect 251652 381942 251712 381970
rect 251974 381956 252002 382214
rect 252112 381970 252140 385222
rect 252480 381970 252508 388554
rect 252664 385286 252692 589902
rect 252928 393372 252980 393378
rect 252928 393314 252980 393320
rect 252744 391400 252796 391406
rect 252744 391342 252796 391348
rect 252652 385280 252704 385286
rect 252652 385222 252704 385228
rect 252756 381970 252784 391342
rect 252940 385150 252968 393314
rect 253020 392828 253072 392834
rect 253020 392770 253072 392776
rect 252928 385144 252980 385150
rect 252928 385086 252980 385092
rect 253032 381970 253060 392770
rect 253216 390590 253244 683130
rect 254032 399764 254084 399770
rect 254032 399706 254084 399712
rect 253480 391468 253532 391474
rect 253480 391410 253532 391416
rect 253204 390584 253256 390590
rect 253204 390526 253256 390532
rect 253204 385280 253256 385286
rect 253204 385222 253256 385228
rect 253216 381970 253244 385222
rect 253492 381970 253520 391410
rect 253848 385348 253900 385354
rect 253848 385290 253900 385296
rect 253860 385150 253888 385290
rect 254044 385218 254072 399706
rect 254584 394188 254636 394194
rect 254584 394130 254636 394136
rect 254400 391536 254452 391542
rect 254400 391478 254452 391484
rect 254308 388748 254360 388754
rect 254308 388690 254360 388696
rect 254032 385212 254084 385218
rect 254032 385154 254084 385160
rect 253756 385144 253808 385150
rect 253756 385086 253808 385092
rect 253848 385144 253900 385150
rect 253848 385086 253900 385092
rect 253768 381970 253796 385086
rect 254320 381970 254348 388690
rect 252112 381942 252264 381970
rect 252480 381942 252540 381970
rect 252756 381942 252816 381970
rect 252928 381948 252980 381954
rect 253032 381942 253092 381970
rect 253216 381942 253368 381970
rect 253492 381942 253644 381970
rect 253768 381942 253920 381970
rect 254196 381942 254348 381970
rect 254412 381970 254440 391478
rect 254596 381970 254624 394130
rect 254952 388884 255004 388890
rect 254952 388826 255004 388832
rect 254412 381942 254472 381970
rect 254596 381942 254748 381970
rect 252928 381890 252980 381896
rect 249168 381806 249228 381834
rect 250720 381744 250772 381750
rect 250720 381686 250772 381692
rect 250732 381546 250760 381686
rect 252940 381614 252968 381890
rect 254964 381834 254992 388826
rect 255136 385212 255188 385218
rect 255136 385154 255188 385160
rect 255148 381970 255176 385154
rect 255608 382242 255636 700470
rect 265624 700460 265676 700466
rect 265624 700402 265676 700408
rect 257620 700392 257672 700398
rect 257620 700334 257672 700340
rect 257344 683256 257396 683262
rect 257344 683198 257396 683204
rect 256792 590096 256844 590102
rect 256792 590038 256844 590044
rect 256240 392896 256292 392902
rect 256240 392838 256292 392844
rect 255964 388816 256016 388822
rect 255964 388758 256016 388764
rect 255688 387456 255740 387462
rect 255688 387398 255740 387404
rect 255562 382214 255636 382242
rect 255148 381942 255300 381970
rect 255562 381956 255590 382214
rect 255700 381970 255728 387398
rect 255976 381970 256004 388758
rect 256252 381970 256280 392838
rect 256516 387388 256568 387394
rect 256516 387330 256568 387336
rect 256528 381970 256556 387330
rect 256804 381970 256832 590038
rect 257160 394120 257212 394126
rect 257160 394062 257212 394068
rect 257068 382016 257120 382022
rect 255700 381942 255852 381970
rect 255976 381942 256128 381970
rect 256252 381942 256404 381970
rect 256528 381942 256680 381970
rect 256804 381942 256956 381970
rect 257068 381958 257120 381964
rect 257172 381970 257200 394062
rect 257356 386510 257384 683198
rect 257436 590028 257488 590034
rect 257436 589970 257488 589976
rect 257344 386504 257396 386510
rect 257344 386446 257396 386452
rect 257448 381970 257476 589970
rect 257632 402974 257660 700334
rect 258724 700324 258776 700330
rect 258724 700266 258776 700272
rect 257632 402946 257936 402974
rect 257620 389972 257672 389978
rect 257620 389914 257672 389920
rect 257632 381970 257660 389914
rect 257908 381970 257936 402946
rect 258736 393378 258764 700266
rect 264244 696992 264296 696998
rect 264244 696934 264296 696940
rect 258816 670812 258868 670818
rect 258816 670754 258868 670760
rect 258724 393372 258776 393378
rect 258724 393314 258776 393320
rect 258724 392012 258776 392018
rect 258724 391954 258776 391960
rect 258540 391332 258592 391338
rect 258540 391274 258592 391280
rect 258172 388680 258224 388686
rect 258172 388622 258224 388628
rect 258184 381970 258212 388622
rect 258552 381970 258580 391274
rect 258632 382968 258684 382974
rect 258632 382910 258684 382916
rect 258644 382634 258672 382910
rect 258632 382628 258684 382634
rect 258632 382570 258684 382576
rect 258736 381970 258764 391954
rect 258828 390590 258856 670754
rect 261484 643136 261536 643142
rect 261484 643078 261536 643084
rect 259828 632120 259880 632126
rect 259828 632062 259880 632068
rect 259552 605872 259604 605878
rect 259552 605814 259604 605820
rect 259276 391604 259328 391610
rect 259276 391546 259328 391552
rect 258816 390584 258868 390590
rect 258816 390526 258868 390532
rect 259000 386504 259052 386510
rect 259000 386446 259052 386452
rect 259012 381970 259040 386446
rect 259288 381970 259316 391546
rect 259564 385218 259592 605814
rect 259552 385212 259604 385218
rect 259552 385154 259604 385160
rect 259642 383616 259698 383625
rect 259642 383551 259698 383560
rect 259656 382945 259684 383551
rect 259642 382936 259698 382945
rect 259642 382871 259698 382880
rect 259656 381970 259684 382871
rect 259840 381970 259868 632062
rect 260472 393440 260524 393446
rect 260472 393382 260524 393388
rect 260196 390584 260248 390590
rect 260196 390526 260248 390532
rect 260104 385212 260156 385218
rect 260104 385154 260156 385160
rect 260116 381970 260144 385154
rect 260208 383625 260236 390526
rect 260194 383616 260250 383625
rect 260194 383551 260250 383560
rect 260484 381970 260512 393382
rect 260932 391264 260984 391270
rect 260932 391206 260984 391212
rect 260656 387252 260708 387258
rect 260656 387194 260708 387200
rect 260668 381970 260696 387194
rect 260944 381970 260972 391206
rect 261496 390182 261524 643078
rect 261576 590708 261628 590714
rect 261576 590650 261628 590656
rect 261484 390176 261536 390182
rect 261484 390118 261536 390124
rect 261588 390114 261616 590650
rect 261668 474768 261720 474774
rect 261668 474710 261720 474716
rect 261576 390108 261628 390114
rect 261576 390050 261628 390056
rect 261300 388544 261352 388550
rect 261300 388486 261352 388492
rect 261208 383852 261260 383858
rect 261208 383794 261260 383800
rect 254964 381806 255024 381834
rect 256240 381812 256292 381818
rect 256240 381754 256292 381760
rect 255136 381744 255188 381750
rect 255136 381686 255188 381692
rect 252928 381608 252980 381614
rect 252928 381550 252980 381556
rect 250720 381540 250772 381546
rect 250720 381482 250772 381488
rect 255148 381478 255176 381686
rect 256252 381478 256280 381754
rect 257080 381478 257108 381958
rect 257172 381942 257232 381970
rect 257448 381942 257508 381970
rect 257632 381942 257784 381970
rect 257908 381942 258060 381970
rect 258184 381942 258336 381970
rect 258552 381942 258612 381970
rect 258736 381942 258888 381970
rect 259012 381942 259164 381970
rect 259288 381942 259440 381970
rect 259656 381942 259716 381970
rect 259840 381942 259992 381970
rect 260116 381942 260268 381970
rect 260484 381942 260544 381970
rect 260668 381942 260820 381970
rect 260944 381942 261096 381970
rect 257908 381857 257936 381942
rect 257894 381848 257950 381857
rect 257894 381783 257950 381792
rect 259828 381744 259880 381750
rect 259828 381686 259880 381692
rect 259840 381478 259868 381686
rect 261220 381682 261248 383794
rect 261312 383722 261340 388486
rect 261484 388476 261536 388482
rect 261484 388418 261536 388424
rect 261300 383716 261352 383722
rect 261300 383658 261352 383664
rect 261312 381970 261340 383658
rect 261496 381970 261524 388418
rect 261680 386510 261708 474710
rect 262588 448588 262640 448594
rect 262588 448530 262640 448536
rect 261760 422340 261812 422346
rect 261760 422282 261812 422288
rect 261772 386578 261800 422282
rect 262128 393984 262180 393990
rect 262128 393926 262180 393932
rect 261944 392760 261996 392766
rect 261944 392702 261996 392708
rect 261760 386572 261812 386578
rect 261760 386514 261812 386520
rect 261668 386504 261720 386510
rect 261668 386446 261720 386452
rect 261956 382242 261984 392702
rect 262140 384305 262168 393926
rect 262312 386504 262364 386510
rect 262312 386446 262364 386452
rect 262126 384296 262182 384305
rect 262126 384231 262182 384240
rect 261910 382214 261984 382242
rect 261312 381942 261372 381970
rect 261496 381942 261648 381970
rect 261910 381956 261938 382214
rect 262140 381970 262168 384231
rect 262324 381970 262352 386446
rect 262600 381970 262628 448530
rect 263784 409896 263836 409902
rect 263784 409838 263836 409844
rect 263416 397520 263468 397526
rect 263416 397462 263468 397468
rect 263140 386572 263192 386578
rect 263140 386514 263192 386520
rect 262864 385280 262916 385286
rect 262864 385222 262916 385228
rect 262876 381970 262904 385222
rect 263152 381970 263180 386514
rect 263428 381970 263456 397462
rect 263796 381970 263824 409838
rect 264256 390046 264284 696934
rect 265636 394194 265664 700402
rect 267660 697610 267688 703520
rect 283852 700534 283880 703520
rect 283840 700528 283892 700534
rect 283840 700470 283892 700476
rect 266360 697604 266412 697610
rect 266360 697546 266412 697552
rect 267648 697604 267700 697610
rect 267648 697546 267700 697552
rect 266372 399770 266400 697546
rect 279424 536852 279476 536858
rect 279424 536794 279476 536800
rect 278044 535492 278096 535498
rect 278044 535434 278096 535440
rect 275284 532772 275336 532778
rect 275284 532714 275336 532720
rect 273904 529984 273956 529990
rect 273904 529926 273956 529932
rect 271144 507884 271196 507890
rect 271144 507826 271196 507832
rect 266360 399764 266412 399770
rect 266360 399706 266412 399712
rect 265624 394188 265676 394194
rect 265624 394130 265676 394136
rect 264244 390040 264296 390046
rect 264244 389982 264296 389988
rect 271156 389174 271184 507826
rect 273916 395962 273944 529926
rect 273996 528624 274048 528630
rect 273996 528566 274048 528572
rect 274008 396030 274036 528566
rect 275296 397390 275324 532714
rect 277308 398132 277360 398138
rect 277308 398074 277360 398080
rect 275284 397384 275336 397390
rect 275284 397326 275336 397332
rect 273996 396024 274048 396030
rect 273996 395966 274048 395972
rect 273904 395956 273956 395962
rect 273904 395898 273956 395904
rect 271972 395412 272024 395418
rect 271972 395354 272024 395360
rect 271984 390046 272012 395354
rect 272524 395344 272576 395350
rect 272524 395286 272576 395292
rect 271972 390040 272024 390046
rect 271972 389982 272024 389988
rect 271156 389146 271552 389174
rect 271524 386374 271552 389146
rect 271512 386368 271564 386374
rect 271512 386310 271564 386316
rect 270866 385112 270922 385121
rect 270866 385047 270922 385056
rect 267004 384804 267056 384810
rect 267004 384746 267056 384752
rect 264888 384328 264940 384334
rect 264888 384270 264940 384276
rect 264520 383920 264572 383926
rect 264520 383862 264572 383868
rect 264060 382968 264112 382974
rect 264060 382910 264112 382916
rect 263968 382016 264020 382022
rect 262140 381942 262200 381970
rect 262324 381942 262476 381970
rect 262600 381942 262752 381970
rect 262876 381942 263028 381970
rect 263152 381942 263304 381970
rect 263428 381942 263580 381970
rect 263796 381942 263856 381970
rect 263968 381958 264020 381964
rect 261208 381676 261260 381682
rect 261208 381618 261260 381624
rect 263980 381478 264008 381958
rect 264072 381834 264100 382910
rect 264244 382900 264296 382906
rect 264244 382842 264296 382848
rect 264256 381970 264284 382842
rect 264532 381970 264560 383862
rect 264796 383036 264848 383042
rect 264796 382978 264848 382984
rect 264808 381970 264836 382978
rect 264900 382974 264928 384270
rect 266450 384160 266506 384169
rect 266450 384095 266506 384104
rect 264888 382968 264940 382974
rect 264888 382910 264940 382916
rect 266176 382492 266228 382498
rect 266176 382434 266228 382440
rect 265348 382424 265400 382430
rect 265348 382366 265400 382372
rect 265072 382356 265124 382362
rect 265072 382298 265124 382304
rect 265084 381970 265112 382298
rect 265360 381970 265388 382366
rect 265624 382288 265676 382294
rect 265624 382230 265676 382236
rect 265636 381970 265664 382230
rect 265900 382016 265952 382022
rect 264256 381942 264408 381970
rect 264532 381942 264684 381970
rect 264808 381942 264960 381970
rect 265084 381942 265236 381970
rect 265360 381942 265512 381970
rect 265636 381942 265788 381970
rect 266188 381970 266216 382434
rect 266464 381970 266492 384095
rect 267016 381970 267044 384746
rect 270316 384668 270368 384674
rect 270316 384610 270368 384616
rect 267648 384464 267700 384470
rect 267646 384432 267648 384441
rect 267700 384432 267702 384441
rect 267646 384367 267702 384376
rect 268198 384432 268254 384441
rect 268198 384367 268254 384376
rect 269764 384396 269816 384402
rect 267554 382800 267610 382809
rect 267554 382735 267610 382744
rect 267568 381970 267596 382735
rect 267832 382560 267884 382566
rect 267832 382502 267884 382508
rect 267844 381970 267872 382502
rect 268212 381970 268240 384367
rect 269764 384338 269816 384344
rect 269488 384260 269540 384266
rect 269488 384202 269540 384208
rect 268658 384024 268714 384033
rect 268658 383959 268714 383968
rect 268382 382664 268438 382673
rect 268382 382599 268438 382608
rect 268396 381970 268424 382599
rect 268672 381970 268700 383959
rect 269500 381970 269528 384202
rect 269776 381970 269804 384338
rect 270040 383784 270092 383790
rect 270040 383726 270092 383732
rect 270052 381970 270080 383726
rect 270328 381970 270356 384610
rect 270880 381970 270908 385047
rect 271418 383344 271474 383353
rect 271418 383279 271474 383288
rect 271432 381970 271460 383279
rect 265952 381964 266064 381970
rect 265900 381958 266064 381964
rect 265912 381942 266064 381958
rect 266188 381942 266340 381970
rect 266464 381942 266616 381970
rect 267016 381942 267168 381970
rect 267292 381954 267444 381970
rect 267280 381948 267444 381954
rect 267332 381942 267444 381948
rect 267568 381942 267720 381970
rect 267844 381942 267996 381970
rect 268212 381942 268272 381970
rect 268396 381942 268548 381970
rect 268672 381942 268824 381970
rect 269500 381942 269652 381970
rect 269776 381942 269928 381970
rect 270052 381942 270204 381970
rect 270328 381942 270480 381970
rect 270880 381942 271032 381970
rect 271308 381942 271460 381970
rect 271524 381970 271552 386310
rect 272536 386306 272564 395286
rect 272616 394052 272668 394058
rect 272616 393994 272668 394000
rect 272524 386300 272576 386306
rect 272524 386242 272576 386248
rect 272628 386238 272656 393994
rect 274008 393314 274036 395966
rect 274180 395956 274232 395962
rect 274180 395898 274232 395904
rect 273640 393286 274036 393314
rect 273076 390516 273128 390522
rect 273076 390458 273128 390464
rect 273088 390046 273116 390458
rect 273076 390040 273128 390046
rect 273076 389982 273128 389988
rect 273088 389174 273116 389982
rect 273088 389146 273208 389174
rect 272800 386300 272852 386306
rect 272800 386242 272852 386248
rect 272248 386232 272300 386238
rect 272248 386174 272300 386180
rect 272616 386232 272668 386238
rect 272616 386174 272668 386180
rect 272260 381970 272288 386174
rect 272524 382492 272576 382498
rect 272524 382434 272576 382440
rect 272536 381970 272564 382434
rect 272812 381970 272840 386242
rect 273074 384704 273130 384713
rect 273074 384639 273130 384648
rect 273088 381970 273116 384639
rect 271524 381942 271584 381970
rect 272136 381942 272288 381970
rect 272412 381942 272564 381970
rect 272688 381942 272840 381970
rect 272964 381942 273116 381970
rect 273180 381970 273208 389146
rect 273442 384840 273498 384849
rect 273442 384775 273498 384784
rect 273456 381970 273484 384775
rect 273640 381970 273668 393286
rect 274192 381970 274220 395898
rect 274824 385756 274876 385762
rect 274824 385698 274876 385704
rect 274456 384192 274508 384198
rect 274456 384134 274508 384140
rect 274468 381970 274496 384134
rect 274548 383716 274600 383722
rect 274548 383658 274600 383664
rect 274560 382129 274588 383658
rect 274546 382120 274602 382129
rect 274546 382055 274602 382064
rect 273180 381942 273240 381970
rect 273456 381942 273516 381970
rect 273640 381942 273792 381970
rect 274192 381942 274344 381970
rect 274468 381942 274620 381970
rect 267280 381890 267332 381896
rect 268936 381880 268988 381886
rect 264072 381806 264132 381834
rect 269210 381848 269266 381857
rect 268988 381828 269100 381834
rect 268936 381822 269100 381828
rect 268948 381806 269100 381822
rect 273902 381848 273958 381857
rect 269266 381806 269376 381834
rect 269210 381783 269266 381792
rect 274836 381834 274864 385698
rect 275008 382832 275060 382838
rect 275008 382774 275060 382780
rect 275020 381970 275048 382774
rect 275296 381970 275324 397326
rect 275928 396772 275980 396778
rect 275928 396714 275980 396720
rect 275940 396098 275968 396714
rect 275376 396092 275428 396098
rect 275376 396034 275428 396040
rect 275928 396092 275980 396098
rect 275928 396034 275980 396040
rect 275388 386442 275416 396034
rect 277320 395962 277348 398074
rect 277308 395956 277360 395962
rect 277308 395898 277360 395904
rect 277320 393314 277348 395898
rect 276952 393286 277348 393314
rect 275376 386436 275428 386442
rect 275376 386378 275428 386384
rect 275836 386436 275888 386442
rect 275836 386378 275888 386384
rect 275560 383988 275612 383994
rect 275560 383930 275612 383936
rect 275572 381970 275600 383930
rect 275848 381970 275876 386378
rect 276480 385688 276532 385694
rect 276480 385630 276532 385636
rect 276492 381970 276520 385630
rect 276754 382528 276810 382537
rect 276754 382463 276810 382472
rect 276768 381970 276796 382463
rect 276952 381970 276980 393286
rect 278056 385694 278084 535434
rect 278136 534132 278188 534138
rect 278136 534074 278188 534080
rect 278148 396098 278176 534074
rect 278228 531344 278280 531350
rect 278228 531286 278280 531292
rect 278136 396092 278188 396098
rect 278136 396034 278188 396040
rect 278136 385824 278188 385830
rect 278136 385766 278188 385772
rect 278044 385688 278096 385694
rect 278044 385630 278096 385636
rect 278042 382664 278098 382673
rect 278042 382599 278098 382608
rect 278056 381970 278084 382599
rect 275020 381942 275172 381970
rect 275296 381942 275448 381970
rect 275572 381942 275724 381970
rect 275848 381942 276000 381970
rect 276492 381942 276552 381970
rect 276768 381942 276828 381970
rect 276952 381942 277104 381970
rect 277932 381942 278084 381970
rect 278148 381970 278176 385766
rect 278240 385762 278268 531286
rect 278596 399560 278648 399566
rect 278596 399502 278648 399508
rect 278228 385756 278280 385762
rect 278228 385698 278280 385704
rect 278410 382392 278466 382401
rect 278410 382327 278466 382336
rect 278424 381970 278452 382327
rect 278608 381970 278636 399502
rect 279148 396840 279200 396846
rect 279148 396782 279200 396788
rect 278964 382832 279016 382838
rect 278964 382774 279016 382780
rect 278976 381970 279004 382774
rect 279160 381970 279188 396782
rect 279436 395962 279464 536794
rect 295984 509312 296036 509318
rect 295984 509254 296036 509260
rect 287428 497208 287480 497214
rect 287428 497150 287480 497156
rect 279700 497072 279752 497078
rect 279700 497014 279752 497020
rect 279424 395956 279476 395962
rect 279424 395898 279476 395904
rect 279516 384260 279568 384266
rect 279516 384202 279568 384208
rect 279528 381970 279556 384202
rect 279712 381970 279740 497014
rect 282184 497004 282236 497010
rect 282184 496946 282236 496952
rect 281908 414724 281960 414730
rect 281908 414666 281960 414672
rect 281920 402974 281948 414666
rect 281920 402946 282132 402974
rect 281816 400988 281868 400994
rect 281816 400930 281868 400936
rect 280252 399628 280304 399634
rect 280252 399570 280304 399576
rect 280264 385218 280292 399570
rect 280804 399492 280856 399498
rect 280804 399434 280856 399440
rect 280344 398200 280396 398206
rect 280344 398142 280396 398148
rect 280252 385212 280304 385218
rect 280252 385154 280304 385160
rect 280068 382288 280120 382294
rect 280068 382230 280120 382236
rect 280080 381970 280108 382230
rect 280356 381970 280384 398142
rect 280528 382764 280580 382770
rect 280528 382706 280580 382712
rect 280540 381970 280568 382706
rect 280816 381970 280844 399434
rect 281828 389174 281856 400930
rect 281828 389146 281948 389174
rect 281632 386504 281684 386510
rect 281632 386446 281684 386452
rect 281356 385212 281408 385218
rect 281356 385154 281408 385160
rect 281078 384568 281134 384577
rect 281078 384503 281134 384512
rect 281092 381970 281120 384503
rect 281368 381970 281396 385154
rect 281644 381970 281672 386446
rect 281920 381970 281948 389146
rect 282104 382106 282132 402946
rect 282196 385014 282224 496946
rect 285220 496936 285272 496942
rect 285220 496878 285272 496884
rect 285772 496936 285824 496942
rect 285772 496878 285824 496884
rect 284392 414860 284444 414866
rect 284392 414802 284444 414808
rect 283656 414792 283708 414798
rect 283656 414734 283708 414740
rect 283012 401056 283064 401062
rect 283012 400998 283064 401004
rect 283024 388482 283052 400998
rect 283104 400920 283156 400926
rect 283104 400862 283156 400868
rect 283012 388476 283064 388482
rect 283012 388418 283064 388424
rect 282184 385008 282236 385014
rect 282184 384950 282236 384956
rect 282104 382078 282500 382106
rect 282472 381970 282500 382078
rect 283116 381970 283144 400862
rect 283564 383716 283616 383722
rect 283564 383658 283616 383664
rect 283576 381970 283604 383658
rect 278148 381942 278208 381970
rect 278424 381942 278484 381970
rect 278608 381942 278760 381970
rect 278976 381942 279036 381970
rect 279160 381942 279312 381970
rect 279528 381942 279588 381970
rect 279712 381942 279864 381970
rect 280080 381942 280140 381970
rect 280356 381942 280416 381970
rect 280540 381942 280692 381970
rect 280816 381942 280968 381970
rect 281092 381942 281244 381970
rect 281368 381942 281520 381970
rect 281644 381942 281796 381970
rect 281920 381942 282072 381970
rect 282472 381942 282624 381970
rect 283116 381942 283176 381970
rect 283452 381942 283604 381970
rect 283668 381970 283696 414734
rect 284404 402974 284432 414802
rect 284404 402946 284708 402974
rect 284116 388476 284168 388482
rect 284116 388418 284168 388424
rect 283976 382120 284032 382129
rect 283976 382055 284032 382064
rect 283668 381942 283728 381970
rect 283990 381956 284018 382055
rect 284128 381970 284156 388418
rect 284484 382628 284536 382634
rect 284484 382570 284536 382576
rect 284496 381970 284524 382570
rect 284680 381970 284708 402946
rect 285128 383920 285180 383926
rect 285128 383862 285180 383868
rect 285140 382242 285168 383862
rect 285094 382214 285168 382242
rect 284128 381942 284280 381970
rect 284496 381942 284556 381970
rect 284680 381942 284832 381970
rect 285094 381956 285122 382214
rect 285232 381970 285260 496878
rect 285784 388482 285812 496878
rect 287152 496868 287204 496874
rect 287152 496810 287204 496816
rect 285864 399696 285916 399702
rect 285864 399638 285916 399644
rect 285772 388476 285824 388482
rect 285772 388418 285824 388424
rect 285588 384668 285640 384674
rect 285588 384610 285640 384616
rect 285600 381970 285628 384610
rect 285876 381970 285904 399638
rect 287164 389774 287192 496810
rect 287152 389768 287204 389774
rect 287152 389710 287204 389716
rect 286876 388476 286928 388482
rect 286876 388418 286928 388424
rect 286324 385008 286376 385014
rect 286324 384950 286376 384956
rect 286140 382560 286192 382566
rect 286140 382502 286192 382508
rect 285232 381942 285384 381970
rect 285600 381942 285660 381970
rect 285876 381942 285936 381970
rect 276110 381848 276166 381857
rect 273958 381806 274068 381834
rect 274836 381806 274896 381834
rect 273902 381783 273958 381792
rect 277766 381848 277822 381857
rect 276166 381806 276276 381834
rect 277656 381806 277766 381834
rect 276110 381783 276166 381792
rect 282458 381848 282514 381857
rect 282348 381806 282458 381834
rect 277766 381783 277822 381792
rect 286152 381834 286180 382502
rect 286336 381970 286364 384950
rect 286784 384804 286836 384810
rect 286784 384746 286836 384752
rect 286796 382242 286824 384746
rect 286750 382214 286824 382242
rect 286336 381942 286488 381970
rect 286750 381956 286778 382214
rect 286888 381970 286916 388418
rect 287244 382356 287296 382362
rect 287244 382298 287296 382304
rect 287256 381970 287284 382298
rect 287440 381970 287468 497150
rect 288624 497140 288676 497146
rect 288624 497082 288676 497088
rect 288532 497072 288584 497078
rect 288532 497014 288584 497020
rect 287980 389768 288032 389774
rect 287980 389710 288032 389716
rect 287886 383752 287942 383761
rect 287886 383687 287942 383696
rect 287900 382242 287928 383687
rect 287854 382214 287928 382242
rect 286888 381942 287040 381970
rect 287256 381942 287316 381970
rect 287440 381942 287592 381970
rect 287854 381956 287882 382214
rect 287992 381970 288020 389710
rect 288544 389366 288572 497014
rect 288532 389360 288584 389366
rect 288532 389302 288584 389308
rect 288530 381984 288586 381993
rect 287992 381942 288144 381970
rect 288420 381942 288530 381970
rect 288636 381970 288664 497082
rect 292672 497004 292724 497010
rect 292672 496946 292724 496952
rect 291292 414724 291344 414730
rect 291292 414666 291344 414672
rect 290740 395412 290792 395418
rect 290740 395354 290792 395360
rect 289636 389360 289688 389366
rect 289636 389302 289688 389308
rect 289268 385688 289320 385694
rect 289268 385630 289320 385636
rect 289084 382424 289136 382430
rect 289084 382366 289136 382372
rect 289096 381970 289124 382366
rect 289280 382242 289308 385630
rect 288636 381942 288696 381970
rect 288972 381942 289124 381970
rect 289234 382214 289308 382242
rect 289234 381956 289262 382214
rect 289358 381984 289414 381993
rect 288530 381919 288586 381928
rect 289648 381970 289676 389302
rect 290188 388408 290240 388414
rect 290188 388350 290240 388356
rect 289728 384124 289780 384130
rect 289728 384066 289780 384072
rect 289740 384033 289768 384066
rect 289726 384024 289782 384033
rect 289726 383959 289782 383968
rect 290002 382120 290058 382129
rect 290002 382055 290058 382064
rect 290016 381970 290044 382055
rect 290200 381970 290228 388350
rect 290648 383852 290700 383858
rect 290648 383794 290700 383800
rect 290660 382242 290688 383794
rect 290614 382214 290688 382242
rect 289414 381942 289524 381970
rect 289648 381942 289800 381970
rect 290016 381942 290076 381970
rect 290200 381942 290352 381970
rect 290614 381956 290642 382214
rect 290752 381970 290780 395354
rect 290922 384160 290978 384169
rect 291304 384130 291332 414666
rect 292684 402974 292712 496946
rect 295616 426420 295668 426426
rect 295616 426362 295668 426368
rect 292684 402946 292896 402974
rect 291384 394120 291436 394126
rect 291384 394062 291436 394068
rect 290922 384095 290978 384104
rect 291292 384124 291344 384130
rect 290936 384062 290964 384095
rect 291292 384066 291344 384072
rect 290924 384056 290976 384062
rect 290924 383998 290976 384004
rect 291108 383716 291160 383722
rect 291108 383658 291160 383664
rect 291120 382974 291148 383658
rect 291108 382968 291160 382974
rect 291108 382910 291160 382916
rect 291106 382800 291162 382809
rect 291106 382735 291162 382744
rect 291120 381970 291148 382735
rect 291396 381970 291424 394062
rect 292396 394052 292448 394058
rect 292396 393994 292448 394000
rect 291844 384464 291896 384470
rect 291842 384432 291844 384441
rect 291896 384432 291898 384441
rect 291842 384367 291898 384376
rect 291844 384124 291896 384130
rect 291844 384066 291896 384072
rect 291752 384056 291804 384062
rect 291752 383998 291804 384004
rect 291764 382242 291792 383998
rect 291718 382214 291792 382242
rect 290752 381942 290904 381970
rect 291120 381942 291180 381970
rect 291396 381942 291456 381970
rect 291718 381956 291746 382214
rect 291856 381970 291884 384066
rect 292118 381984 292174 381993
rect 291856 381942 292008 381970
rect 289358 381919 289414 381928
rect 292408 381970 292436 393994
rect 292764 383784 292816 383790
rect 292764 383726 292816 383732
rect 292776 381970 292804 383726
rect 292868 383654 292896 402946
rect 294052 396772 294104 396778
rect 294052 396714 294104 396720
rect 293500 393984 293552 393990
rect 293500 393926 293552 393932
rect 293408 383988 293460 383994
rect 293408 383930 293460 383936
rect 292868 383626 292988 383654
rect 292960 381970 292988 383626
rect 293420 382242 293448 383930
rect 293374 382214 293448 382242
rect 292174 381942 292284 381970
rect 292408 381942 292560 381970
rect 292776 381942 292836 381970
rect 292960 381942 293112 381970
rect 293374 381956 293402 382214
rect 293512 381970 293540 393926
rect 294064 388482 294092 396714
rect 294144 395480 294196 395486
rect 294144 395422 294196 395428
rect 294052 388476 294104 388482
rect 294052 388418 294104 388424
rect 293776 384736 293828 384742
rect 293776 384678 293828 384684
rect 293512 381942 293664 381970
rect 292118 381919 292174 381928
rect 286152 381806 286212 381834
rect 282458 381783 282514 381792
rect 270592 381744 270644 381750
rect 270644 381692 270756 381698
rect 270592 381686 270756 381692
rect 270604 381670 270756 381686
rect 276940 381676 276992 381682
rect 276940 381618 276992 381624
rect 282184 381676 282236 381682
rect 282184 381618 282236 381624
rect 276952 381478 276980 381618
rect 277380 381546 277532 381562
rect 277380 381540 277544 381546
rect 277380 381534 277492 381540
rect 277492 381482 277544 381488
rect 282196 381478 282224 381618
rect 293788 381614 293816 384678
rect 293912 382120 293968 382129
rect 293912 382055 293968 382064
rect 293926 381956 293954 382055
rect 294156 381970 294184 395422
rect 294604 395344 294656 395350
rect 294604 395286 294656 395292
rect 294512 383716 294564 383722
rect 294512 383658 294564 383664
rect 294524 382242 294552 383658
rect 294478 382214 294552 382242
rect 294156 381942 294216 381970
rect 294478 381956 294506 382214
rect 294616 381970 294644 395286
rect 295156 388476 295208 388482
rect 295156 388418 295208 388424
rect 294878 381984 294934 381993
rect 294616 381942 294768 381970
rect 295168 381970 295196 388418
rect 295628 384985 295656 426362
rect 295996 397458 296024 509254
rect 296076 507952 296128 507958
rect 296076 507894 296128 507900
rect 296088 426426 296116 507894
rect 296076 426420 296128 426426
rect 296076 426362 296128 426368
rect 295984 397452 296036 397458
rect 295984 397394 296036 397400
rect 295996 393314 296024 397394
rect 295812 393286 296024 393314
rect 295614 384976 295670 384985
rect 295614 384911 295670 384920
rect 295340 384872 295392 384878
rect 295338 384840 295340 384849
rect 295392 384840 295394 384849
rect 295338 384775 295394 384784
rect 295706 381984 295762 381993
rect 294934 381942 295044 381970
rect 295168 381942 295320 381970
rect 295596 381942 295706 381970
rect 294878 381919 294934 381928
rect 295812 381970 295840 393286
rect 299492 388890 299520 703582
rect 299952 703474 299980 703582
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429212 703582 429700 703610
rect 300136 703474 300164 703520
rect 299952 703446 300164 703474
rect 331864 700528 331916 700534
rect 331864 700470 331916 700476
rect 324964 700392 325016 700398
rect 324964 700334 325016 700340
rect 324976 391542 325004 700334
rect 324964 391536 325016 391542
rect 324964 391478 325016 391484
rect 331876 391474 331904 700470
rect 332520 700398 332548 703520
rect 348804 700466 348832 703520
rect 364996 702434 365024 703520
rect 364352 702406 365024 702434
rect 348792 700460 348844 700466
rect 348792 700402 348844 700408
rect 332508 700392 332560 700398
rect 332508 700334 332560 700340
rect 347044 700392 347096 700398
rect 347044 700334 347096 700340
rect 331864 391468 331916 391474
rect 331864 391410 331916 391416
rect 347056 391406 347084 700334
rect 347044 391400 347096 391406
rect 347044 391342 347096 391348
rect 299480 388884 299532 388890
rect 299480 388826 299532 388832
rect 364352 388754 364380 702406
rect 397472 700534 397500 703520
rect 397460 700528 397512 700534
rect 397460 700470 397512 700476
rect 413664 700330 413692 703520
rect 413652 700324 413704 700330
rect 413652 700266 413704 700272
rect 429212 589966 429240 703582
rect 429672 703474 429700 703582
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494072 703582 494652 703610
rect 429856 703474 429884 703520
rect 429672 703446 429884 703474
rect 462332 700398 462360 703520
rect 478524 702434 478552 703520
rect 477512 702406 478552 702434
rect 462320 700392 462372 700398
rect 462320 700334 462372 700340
rect 429200 589960 429252 589966
rect 429200 589902 429252 589908
rect 376942 537024 376998 537033
rect 376942 536959 376998 536968
rect 376956 536858 376984 536959
rect 376944 536852 376996 536858
rect 376944 536794 376996 536800
rect 377034 535936 377090 535945
rect 377034 535871 377090 535880
rect 377048 535498 377076 535871
rect 377036 535492 377088 535498
rect 377036 535434 377088 535440
rect 376942 534304 376998 534313
rect 376942 534239 376998 534248
rect 376956 534138 376984 534239
rect 376944 534132 376996 534138
rect 376944 534074 376996 534080
rect 377034 533216 377090 533225
rect 377034 533151 377090 533160
rect 377048 532778 377076 533151
rect 377036 532772 377088 532778
rect 377036 532714 377088 532720
rect 376942 531584 376998 531593
rect 376942 531519 376998 531528
rect 376956 531350 376984 531519
rect 376944 531344 376996 531350
rect 376944 531286 376996 531292
rect 376942 530224 376998 530233
rect 376942 530159 376998 530168
rect 376956 529990 376984 530159
rect 376944 529984 376996 529990
rect 376944 529926 376996 529932
rect 376852 528624 376904 528630
rect 376850 528592 376852 528601
rect 376904 528592 376906 528601
rect 376850 528527 376906 528536
rect 471244 510672 471296 510678
rect 471244 510614 471296 510620
rect 376942 510232 376998 510241
rect 376942 510167 376998 510176
rect 376956 509318 376984 510167
rect 376944 509312 376996 509318
rect 376944 509254 376996 509260
rect 377034 508600 377090 508609
rect 377034 508535 377090 508544
rect 376758 508328 376814 508337
rect 376758 508263 376814 508272
rect 376772 507958 376800 508263
rect 376760 507952 376812 507958
rect 376760 507894 376812 507900
rect 377048 507890 377076 508535
rect 377036 507884 377088 507890
rect 377036 507826 377088 507832
rect 397458 498128 397514 498137
rect 397458 498063 397514 498072
rect 425058 498128 425114 498137
rect 425058 498063 425114 498072
rect 397472 497214 397500 498063
rect 409878 497720 409934 497729
rect 409878 497655 409934 497664
rect 398930 497312 398986 497321
rect 398930 497247 398986 497256
rect 403162 497312 403218 497321
rect 403162 497247 403218 497256
rect 397460 497208 397512 497214
rect 397460 497150 397512 497156
rect 398838 497176 398894 497185
rect 398838 497111 398840 497120
rect 398892 497111 398894 497120
rect 398840 497082 398892 497088
rect 398944 497078 398972 497247
rect 398932 497072 398984 497078
rect 398932 497014 398984 497020
rect 403176 497010 403204 497247
rect 404358 497040 404414 497049
rect 403164 497004 403216 497010
rect 404358 496975 404414 496984
rect 403164 496946 403216 496952
rect 404372 496942 404400 496975
rect 404360 496936 404412 496942
rect 391938 496904 391994 496913
rect 391938 496839 391994 496848
rect 393318 496904 393374 496913
rect 393318 496839 393374 496848
rect 394698 496904 394754 496913
rect 394698 496839 394754 496848
rect 400218 496904 400274 496913
rect 400218 496839 400274 496848
rect 401598 496904 401654 496913
rect 404360 496878 404412 496884
rect 404450 496904 404506 496913
rect 401598 496839 401654 496848
rect 404450 496839 404506 496848
rect 405738 496904 405794 496913
rect 409892 496874 409920 497655
rect 415398 496904 415454 496913
rect 405738 496839 405794 496848
rect 409880 496868 409932 496874
rect 364340 388748 364392 388754
rect 364340 388690 364392 388696
rect 391952 386306 391980 496839
rect 393332 386374 393360 496839
rect 394712 390522 394740 496839
rect 400232 395418 400260 496839
rect 401612 414730 401640 496839
rect 401600 414724 401652 414730
rect 401600 414666 401652 414672
rect 404464 395486 404492 496839
rect 405752 396778 405780 496839
rect 415398 496839 415454 496848
rect 419538 496904 419594 496913
rect 419538 496839 419594 496848
rect 409880 496810 409932 496816
rect 405740 396772 405792 396778
rect 405740 396714 405792 396720
rect 404452 395480 404504 395486
rect 404452 395422 404504 395428
rect 400220 395412 400272 395418
rect 400220 395354 400272 395360
rect 394700 390516 394752 390522
rect 394700 390458 394752 390464
rect 393320 386368 393372 386374
rect 393320 386310 393372 386316
rect 391940 386300 391992 386306
rect 391940 386242 391992 386248
rect 415412 385694 415440 496839
rect 419552 388482 419580 496839
rect 425072 394126 425100 498063
rect 429198 496904 429254 496913
rect 429198 496839 429254 496848
rect 434718 496904 434774 496913
rect 434718 496839 434774 496848
rect 440238 496904 440294 496913
rect 440238 496839 440294 496848
rect 425060 394120 425112 394126
rect 425060 394062 425112 394068
rect 429212 394058 429240 496839
rect 429200 394052 429252 394058
rect 429200 393994 429252 394000
rect 434732 393990 434760 496839
rect 440252 395350 440280 496839
rect 440240 395344 440292 395350
rect 440240 395286 440292 395292
rect 434720 393984 434772 393990
rect 434720 393926 434772 393932
rect 419540 388476 419592 388482
rect 419540 388418 419592 388424
rect 471256 387326 471284 510614
rect 477512 392834 477540 702406
rect 477500 392828 477552 392834
rect 477500 392770 477552 392776
rect 494072 388618 494100 703582
rect 494624 703474 494652 703582
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 494808 703474 494836 703520
rect 494624 703446 494836 703474
rect 527192 389910 527220 703520
rect 543476 702434 543504 703520
rect 559668 702434 559696 703520
rect 542372 702406 543504 702434
rect 558932 702406 559696 702434
rect 542372 392698 542400 702406
rect 542360 392692 542412 392698
rect 542360 392634 542412 392640
rect 527180 389904 527232 389910
rect 527180 389846 527232 389852
rect 494060 388612 494112 388618
rect 494060 388554 494112 388560
rect 471244 387320 471296 387326
rect 471244 387262 471296 387268
rect 558932 387190 558960 702406
rect 580170 697232 580226 697241
rect 580170 697167 580226 697176
rect 580184 696998 580212 697167
rect 580172 696992 580224 696998
rect 580172 696934 580224 696940
rect 580170 683904 580226 683913
rect 580170 683839 580226 683848
rect 580184 683194 580212 683839
rect 580172 683188 580224 683194
rect 580172 683130 580224 683136
rect 580172 670744 580224 670750
rect 580170 670712 580172 670721
rect 580224 670712 580226 670721
rect 580170 670647 580226 670656
rect 580170 644056 580226 644065
rect 580170 643991 580226 644000
rect 580184 643142 580212 643991
rect 580172 643136 580224 643142
rect 580172 643078 580224 643084
rect 580170 630864 580226 630873
rect 580170 630799 580226 630808
rect 580184 630698 580212 630799
rect 580172 630692 580224 630698
rect 580172 630634 580224 630640
rect 580170 617536 580226 617545
rect 580170 617471 580226 617480
rect 580184 616894 580212 617471
rect 580172 616888 580224 616894
rect 580172 616830 580224 616836
rect 579802 591016 579858 591025
rect 579802 590951 579858 590960
rect 579816 590714 579844 590951
rect 579804 590708 579856 590714
rect 579804 590650 579856 590656
rect 580354 577688 580410 577697
rect 580354 577623 580410 577632
rect 580262 564360 580318 564369
rect 580262 564295 580318 564304
rect 579618 511320 579674 511329
rect 579618 511255 579674 511264
rect 579632 510678 579660 511255
rect 579620 510672 579672 510678
rect 579620 510614 579672 510620
rect 580170 484664 580226 484673
rect 580170 484599 580226 484608
rect 580184 484430 580212 484599
rect 580172 484424 580224 484430
rect 580172 484366 580224 484372
rect 579986 471472 580042 471481
rect 579986 471407 580042 471416
rect 580000 470626 580028 471407
rect 579988 470620 580040 470626
rect 579988 470562 580040 470568
rect 580170 458144 580226 458153
rect 580170 458079 580226 458088
rect 580184 456822 580212 458079
rect 580172 456816 580224 456822
rect 580172 456758 580224 456764
rect 579618 431624 579674 431633
rect 579618 431559 579674 431568
rect 579632 430642 579660 431559
rect 579620 430636 579672 430642
rect 579620 430578 579672 430584
rect 579710 418296 579766 418305
rect 579710 418231 579766 418240
rect 579724 418198 579752 418231
rect 579712 418192 579764 418198
rect 579712 418134 579764 418140
rect 579986 404968 580042 404977
rect 579986 404903 580042 404912
rect 580000 404394 580028 404903
rect 579988 404388 580040 404394
rect 579988 404330 580040 404336
rect 558920 387184 558972 387190
rect 558920 387126 558972 387132
rect 580276 387122 580304 564295
rect 580368 406434 580396 577623
rect 580446 537840 580502 537849
rect 580446 537775 580502 537784
rect 580356 406428 580408 406434
rect 580356 406370 580408 406376
rect 580460 389842 580488 537775
rect 580538 524512 580594 524521
rect 580538 524447 580594 524456
rect 580552 392630 580580 524447
rect 580540 392624 580592 392630
rect 580540 392566 580592 392572
rect 580448 389836 580500 389842
rect 580448 389778 580500 389784
rect 580264 387116 580316 387122
rect 580264 387058 580316 387064
rect 415400 385688 415452 385694
rect 415400 385630 415452 385636
rect 577964 385144 578016 385150
rect 577964 385086 578016 385092
rect 577780 385076 577832 385082
rect 577780 385018 577832 385024
rect 295982 384976 296038 384985
rect 295982 384911 296038 384920
rect 295996 381970 296024 384911
rect 296812 384804 296864 384810
rect 296812 384746 296864 384752
rect 296536 384056 296588 384062
rect 296536 383998 296588 384004
rect 296258 381984 296314 381993
rect 295812 381942 295872 381970
rect 295996 381942 296258 381970
rect 295706 381919 295762 381928
rect 296548 381970 296576 383998
rect 296626 383752 296682 383761
rect 296626 383687 296682 383696
rect 296424 381942 296576 381970
rect 296640 381970 296668 383687
rect 296640 381942 296700 381970
rect 296258 381919 296314 381928
rect 296824 381682 296852 384746
rect 301872 384668 301924 384674
rect 301872 384610 301924 384616
rect 301780 384328 301832 384334
rect 301780 384270 301832 384276
rect 300124 384192 300176 384198
rect 300124 384134 300176 384140
rect 299480 382288 299532 382294
rect 299480 382230 299532 382236
rect 296812 381676 296864 381682
rect 296812 381618 296864 381624
rect 293776 381608 293828 381614
rect 293776 381550 293828 381556
rect 247408 381472 247460 381478
rect 244260 381414 244424 381420
rect 245474 381440 245530 381449
rect 244260 381398 244412 381414
rect 242714 381375 242770 381384
rect 246026 381440 246082 381449
rect 245530 381398 245640 381426
rect 245474 381375 245530 381384
rect 247408 381414 247460 381420
rect 248236 381472 248288 381478
rect 248236 381414 248288 381420
rect 255136 381472 255188 381478
rect 255136 381414 255188 381420
rect 256240 381472 256292 381478
rect 256240 381414 256292 381420
rect 257068 381472 257120 381478
rect 257068 381414 257120 381420
rect 259828 381472 259880 381478
rect 259828 381414 259880 381420
rect 263968 381472 264020 381478
rect 263968 381414 264020 381420
rect 266728 381472 266780 381478
rect 271972 381472 272024 381478
rect 266780 381420 266892 381426
rect 266728 381414 266892 381420
rect 266740 381398 266892 381414
rect 271860 381420 271972 381426
rect 271860 381414 272024 381420
rect 276940 381472 276992 381478
rect 276940 381414 276992 381420
rect 282184 381472 282236 381478
rect 283012 381472 283064 381478
rect 282184 381414 282236 381420
rect 282900 381420 283012 381426
rect 282900 381414 283064 381420
rect 271860 381398 272012 381414
rect 282900 381398 283052 381414
rect 246026 381375 246082 381384
rect 244096 338564 244148 338570
rect 244096 338506 244148 338512
rect 242992 338020 243044 338026
rect 242992 337962 243044 337968
rect 243004 337278 243032 337962
rect 242992 337272 243044 337278
rect 242992 337214 243044 337220
rect 241428 336932 241480 336938
rect 241428 336874 241480 336880
rect 240048 336864 240100 336870
rect 240048 336806 240100 336812
rect 237378 328264 237434 328273
rect 237378 328199 237434 328208
rect 235998 159352 236054 159361
rect 235998 159287 236054 159296
rect 235908 71732 235960 71738
rect 235908 71674 235960 71680
rect 236012 16574 236040 159287
rect 237392 16574 237420 328199
rect 237472 214600 237524 214606
rect 237470 214568 237472 214577
rect 237524 214568 237526 214577
rect 237470 214503 237526 214512
rect 239586 161120 239642 161129
rect 239586 161055 239642 161064
rect 238758 158128 238814 158137
rect 238758 158063 238814 158072
rect 238772 16574 238800 158063
rect 236012 16546 236592 16574
rect 237392 16546 237696 16574
rect 238772 16546 239352 16574
rect 235816 11688 235868 11694
rect 235816 11630 235868 11636
rect 234632 6886 234752 6914
rect 233884 3596 233936 3602
rect 233884 3538 233936 3544
rect 234632 480 234660 6886
rect 235828 480 235856 11630
rect 232198 354 232310 480
rect 231872 326 232310 354
rect 232198 -960 232310 326
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236564 354 236592 16546
rect 236982 354 237094 480
rect 236564 326 237094 354
rect 237668 354 237696 16546
rect 239324 480 239352 16546
rect 239600 9314 239628 161055
rect 239956 160948 240008 160954
rect 239956 160890 240008 160896
rect 239680 160880 239732 160886
rect 239680 160822 239732 160828
rect 239862 160848 239918 160857
rect 239692 9654 239720 160822
rect 239772 160812 239824 160818
rect 239862 160783 239918 160792
rect 239772 160754 239824 160760
rect 239680 9648 239732 9654
rect 239680 9590 239732 9596
rect 239784 9518 239812 160754
rect 239772 9512 239824 9518
rect 239772 9454 239824 9460
rect 239588 9308 239640 9314
rect 239588 9250 239640 9256
rect 239876 9178 239904 160783
rect 239968 9450 239996 160890
rect 239956 9444 240008 9450
rect 239956 9386 240008 9392
rect 239864 9172 239916 9178
rect 239864 9114 239916 9120
rect 240060 8906 240088 336806
rect 241150 161392 241206 161401
rect 241150 161327 241206 161336
rect 240140 156868 240192 156874
rect 240140 156810 240192 156816
rect 240048 8900 240100 8906
rect 240048 8842 240100 8848
rect 238086 354 238198 480
rect 237668 326 238198 354
rect 236982 -960 237094 326
rect 238086 -960 238198 326
rect 239282 -960 239394 480
rect 240152 354 240180 156810
rect 241164 8974 241192 161327
rect 241242 161256 241298 161265
rect 241242 161191 241298 161200
rect 241256 9246 241284 161191
rect 241336 161016 241388 161022
rect 241336 160958 241388 160964
rect 241348 9382 241376 160958
rect 241336 9376 241388 9382
rect 241336 9318 241388 9324
rect 241244 9240 241296 9246
rect 241244 9182 241296 9188
rect 241152 8968 241204 8974
rect 241152 8910 241204 8916
rect 241440 6050 241468 336874
rect 242348 336728 242400 336734
rect 242348 336670 242400 336676
rect 242164 335844 242216 335850
rect 242164 335786 242216 335792
rect 241520 333804 241572 333810
rect 241520 333746 241572 333752
rect 241532 16574 241560 333746
rect 242072 161084 242124 161090
rect 242072 161026 242124 161032
rect 241532 16546 241744 16574
rect 241428 6044 241480 6050
rect 241428 5986 241480 5992
rect 241716 480 241744 16546
rect 242084 8838 242112 161026
rect 242072 8832 242124 8838
rect 242072 8774 242124 8780
rect 242176 3670 242204 335786
rect 242256 335164 242308 335170
rect 242256 335106 242308 335112
rect 242164 3664 242216 3670
rect 242164 3606 242216 3612
rect 242268 3534 242296 335106
rect 242360 6186 242388 336670
rect 242440 335980 242492 335986
rect 242440 335922 242492 335928
rect 242452 9042 242480 335922
rect 243728 335912 243780 335918
rect 243728 335854 243780 335860
rect 242530 335472 242586 335481
rect 242530 335407 242586 335416
rect 242544 10674 242572 335407
rect 242900 335232 242952 335238
rect 242900 335174 242952 335180
rect 242624 161424 242676 161430
rect 242624 161366 242676 161372
rect 242532 10668 242584 10674
rect 242532 10610 242584 10616
rect 242440 9036 242492 9042
rect 242440 8978 242492 8984
rect 242636 8770 242664 161366
rect 242716 161220 242768 161226
rect 242716 161162 242768 161168
rect 242624 8764 242676 8770
rect 242624 8706 242676 8712
rect 242348 6180 242400 6186
rect 242348 6122 242400 6128
rect 242728 6118 242756 161162
rect 242808 160676 242860 160682
rect 242808 160618 242860 160624
rect 242716 6112 242768 6118
rect 242716 6054 242768 6060
rect 242820 5982 242848 160618
rect 242808 5976 242860 5982
rect 242808 5918 242860 5924
rect 242256 3528 242308 3534
rect 242256 3470 242308 3476
rect 242912 480 242940 335174
rect 243636 332376 243688 332382
rect 243636 332318 243688 332324
rect 243542 331936 243598 331945
rect 243542 331871 243598 331880
rect 242992 158296 243044 158302
rect 242992 158238 243044 158244
rect 243004 16574 243032 158238
rect 243004 16546 243492 16574
rect 243464 3482 243492 16546
rect 243556 3874 243584 331871
rect 243544 3868 243596 3874
rect 243544 3810 243596 3816
rect 243648 3738 243676 332318
rect 243740 7886 243768 335854
rect 243912 335776 243964 335782
rect 243818 335744 243874 335753
rect 243912 335718 243964 335724
rect 243818 335679 243874 335688
rect 243832 89078 243860 335679
rect 243820 89072 243872 89078
rect 243820 89014 243872 89020
rect 243924 89010 243952 335718
rect 244004 161152 244056 161158
rect 244004 161094 244056 161100
rect 243912 89004 243964 89010
rect 243912 88946 243964 88952
rect 244016 9042 244044 161094
rect 244004 9036 244056 9042
rect 244004 8978 244056 8984
rect 243728 7880 243780 7886
rect 243728 7822 243780 7828
rect 244108 6662 244136 338506
rect 244646 338328 244702 338337
rect 244646 338263 244702 338272
rect 244464 337952 244516 337958
rect 244370 337920 244426 337929
rect 244464 337894 244516 337900
rect 244370 337855 244426 337864
rect 244280 337816 244332 337822
rect 244280 337758 244332 337764
rect 244188 336660 244240 336666
rect 244188 336602 244240 336608
rect 244096 6656 244148 6662
rect 244096 6598 244148 6604
rect 244200 3738 244228 336602
rect 244292 5098 244320 337758
rect 244280 5092 244332 5098
rect 244280 5034 244332 5040
rect 244384 4826 244412 337855
rect 244476 178702 244504 337894
rect 244660 336161 244688 338263
rect 291014 338192 291070 338201
rect 291014 338127 291070 338136
rect 244740 338088 244792 338094
rect 290924 338088 290976 338094
rect 244740 338030 244792 338036
rect 244646 336152 244702 336161
rect 244646 336087 244702 336096
rect 244752 329089 244780 338030
rect 244844 338014 245364 338042
rect 244738 329080 244794 329089
rect 244738 329015 244794 329024
rect 244844 323610 244872 338014
rect 245442 337963 245470 338028
rect 245428 337954 245484 337963
rect 245108 337884 245160 337890
rect 245428 337889 245484 337898
rect 245108 337826 245160 337832
rect 244922 337648 244978 337657
rect 244922 337583 244978 337592
rect 244832 323604 244884 323610
rect 244832 323546 244884 323552
rect 244464 178696 244516 178702
rect 244464 178638 244516 178644
rect 244464 159724 244516 159730
rect 244464 159666 244516 159672
rect 244476 16574 244504 159666
rect 244476 16546 244872 16574
rect 244372 4820 244424 4826
rect 244372 4762 244424 4768
rect 243636 3732 243688 3738
rect 243636 3674 243688 3680
rect 244188 3732 244240 3738
rect 244188 3674 244240 3680
rect 244844 3482 244872 16546
rect 244936 3602 244964 337583
rect 245016 337476 245068 337482
rect 245016 337418 245068 337424
rect 245028 336433 245056 337418
rect 245014 336424 245070 336433
rect 245014 336359 245070 336368
rect 245120 336297 245148 337826
rect 245534 337822 245562 338028
rect 245626 337958 245654 338028
rect 245718 337958 245746 338028
rect 245810 337963 245838 338028
rect 245614 337952 245666 337958
rect 245614 337894 245666 337900
rect 245706 337952 245758 337958
rect 245706 337894 245758 337900
rect 245796 337954 245852 337963
rect 245902 337958 245930 338028
rect 245994 337963 246022 338028
rect 245796 337889 245852 337898
rect 245890 337952 245942 337958
rect 245890 337894 245942 337900
rect 245980 337954 246036 337963
rect 245980 337889 246036 337898
rect 245522 337816 245574 337822
rect 246086 337804 246114 338028
rect 246178 337963 246206 338028
rect 246164 337954 246220 337963
rect 246270 337958 246298 338028
rect 246164 337889 246220 337898
rect 246258 337952 246310 337958
rect 246258 337894 246310 337900
rect 246086 337793 246160 337804
rect 246086 337784 246174 337793
rect 246086 337776 246118 337784
rect 245522 337758 245574 337764
rect 245936 337748 245988 337754
rect 246362 337770 246390 338028
rect 246454 337958 246482 338028
rect 246546 337963 246574 338028
rect 246442 337952 246494 337958
rect 246442 337894 246494 337900
rect 246532 337954 246588 337963
rect 246532 337889 246588 337898
rect 246638 337890 246666 338028
rect 246730 337958 246758 338028
rect 246822 337958 246850 338028
rect 246914 337958 246942 338028
rect 246718 337952 246770 337958
rect 246718 337894 246770 337900
rect 246810 337952 246862 337958
rect 246810 337894 246862 337900
rect 246902 337952 246954 337958
rect 247006 337929 247034 338028
rect 247098 337958 247126 338028
rect 247190 337958 247218 338028
rect 247086 337952 247138 337958
rect 246902 337894 246954 337900
rect 246992 337920 247048 337929
rect 246626 337884 246678 337890
rect 247086 337894 247138 337900
rect 247178 337952 247230 337958
rect 247178 337894 247230 337900
rect 247282 337890 247310 338028
rect 247374 337958 247402 338028
rect 247362 337952 247414 337958
rect 247466 337929 247494 338028
rect 247362 337894 247414 337900
rect 247452 337920 247508 337929
rect 246992 337855 247048 337864
rect 247270 337884 247322 337890
rect 246626 337826 246678 337832
rect 247452 337855 247508 337864
rect 247270 337826 247322 337832
rect 247132 337816 247184 337822
rect 246118 337719 246174 337728
rect 246316 337742 246390 337770
rect 246946 337784 247002 337793
rect 246672 337748 246724 337754
rect 245936 337690 245988 337696
rect 245750 337512 245806 337521
rect 245750 337447 245806 337456
rect 245566 336696 245622 336705
rect 245566 336631 245622 336640
rect 245106 336288 245162 336297
rect 245106 336223 245162 336232
rect 245474 336152 245530 336161
rect 245474 336087 245530 336096
rect 245014 335880 245070 335889
rect 245014 335815 245070 335824
rect 245028 13258 245056 335815
rect 245382 335608 245438 335617
rect 245382 335543 245438 335552
rect 245396 333266 245424 335543
rect 245488 335481 245516 336087
rect 245580 335753 245608 336631
rect 245566 335744 245622 335753
rect 245566 335679 245622 335688
rect 245474 335472 245530 335481
rect 245474 335407 245530 335416
rect 245384 333260 245436 333266
rect 245384 333202 245436 333208
rect 245764 330546 245792 337447
rect 245948 334801 245976 337690
rect 246028 337680 246080 337686
rect 246028 337622 246080 337628
rect 245934 334792 245990 334801
rect 245934 334727 245990 334736
rect 246040 331214 246068 337622
rect 246316 331214 246344 337742
rect 246672 337690 246724 337696
rect 246764 337748 246816 337754
rect 247408 337816 247460 337822
rect 247132 337758 247184 337764
rect 247222 337784 247278 337793
rect 246946 337719 247002 337728
rect 246764 337690 246816 337696
rect 246580 337612 246632 337618
rect 246580 337554 246632 337560
rect 246488 337544 246540 337550
rect 246488 337486 246540 337492
rect 246500 331214 246528 337486
rect 245948 331186 246068 331214
rect 246132 331186 246344 331214
rect 246408 331186 246528 331214
rect 245752 330540 245804 330546
rect 245752 330482 245804 330488
rect 245844 330540 245896 330546
rect 245844 330482 245896 330488
rect 245752 330404 245804 330410
rect 245752 330346 245804 330352
rect 245108 320204 245160 320210
rect 245108 320146 245160 320152
rect 245120 97918 245148 320146
rect 245476 161356 245528 161362
rect 245476 161298 245528 161304
rect 245108 97912 245160 97918
rect 245108 97854 245160 97860
rect 245016 13252 245068 13258
rect 245016 13194 245068 13200
rect 245488 6458 245516 161298
rect 245566 160576 245622 160585
rect 245566 160511 245622 160520
rect 245476 6452 245528 6458
rect 245476 6394 245528 6400
rect 245580 6186 245608 160511
rect 245764 9081 245792 330346
rect 245750 9072 245806 9081
rect 245750 9007 245806 9016
rect 245856 8945 245884 330482
rect 245948 10334 245976 331186
rect 246132 330562 246160 331186
rect 246040 330534 246160 330562
rect 246040 13122 246068 330534
rect 246120 330472 246172 330478
rect 246120 330414 246172 330420
rect 246132 177342 246160 330414
rect 246408 316034 246436 331186
rect 246592 330546 246620 337554
rect 246580 330540 246632 330546
rect 246580 330482 246632 330488
rect 246684 330478 246712 337690
rect 246776 336734 246804 337690
rect 246764 336728 246816 336734
rect 246764 336670 246816 336676
rect 246854 336152 246910 336161
rect 246854 336087 246910 336096
rect 246764 332988 246816 332994
rect 246764 332930 246816 332936
rect 246776 331214 246804 332930
rect 246868 332110 246896 336087
rect 246856 332104 246908 332110
rect 246856 332046 246908 332052
rect 246776 331186 246896 331214
rect 246672 330472 246724 330478
rect 246672 330414 246724 330420
rect 246868 325694 246896 331186
rect 246960 330410 246988 337719
rect 247038 337648 247094 337657
rect 247038 337583 247094 337592
rect 247052 334558 247080 337583
rect 247144 335345 247172 337758
rect 247558 337770 247586 338028
rect 247650 337890 247678 338028
rect 247638 337884 247690 337890
rect 247638 337826 247690 337832
rect 247408 337758 247460 337764
rect 247222 337719 247224 337728
rect 247276 337719 247278 337728
rect 247316 337748 247368 337754
rect 247224 337690 247276 337696
rect 247316 337690 247368 337696
rect 247224 337612 247276 337618
rect 247224 337554 247276 337560
rect 247130 335336 247186 335345
rect 247130 335271 247186 335280
rect 247040 334552 247092 334558
rect 247040 334494 247092 334500
rect 247132 333260 247184 333266
rect 247132 333202 247184 333208
rect 246948 330404 247000 330410
rect 246948 330346 247000 330352
rect 246868 325666 246988 325694
rect 246224 316006 246436 316034
rect 246120 177336 246172 177342
rect 246120 177278 246172 177284
rect 246028 13116 246080 13122
rect 246028 13058 246080 13064
rect 245936 10328 245988 10334
rect 245936 10270 245988 10276
rect 245842 8936 245898 8945
rect 245842 8871 245898 8880
rect 245568 6180 245620 6186
rect 245568 6122 245620 6128
rect 246224 4894 246252 316006
rect 246856 160608 246908 160614
rect 246856 160550 246908 160556
rect 246672 158432 246724 158438
rect 246672 158374 246724 158380
rect 246684 6798 246712 158374
rect 246764 158364 246816 158370
rect 246764 158306 246816 158312
rect 246776 6866 246804 158306
rect 246764 6860 246816 6866
rect 246764 6802 246816 6808
rect 246672 6792 246724 6798
rect 246672 6734 246724 6740
rect 246868 6594 246896 160550
rect 246960 100026 246988 325666
rect 247144 320822 247172 333202
rect 247132 320816 247184 320822
rect 247132 320758 247184 320764
rect 246948 100020 247000 100026
rect 246948 99962 247000 99968
rect 247236 10538 247264 337554
rect 247328 333305 247356 337690
rect 247314 333296 247370 333305
rect 247314 333231 247370 333240
rect 247420 333169 247448 337758
rect 247512 337742 247586 337770
rect 247512 336326 247540 337742
rect 247742 337736 247770 338028
rect 247834 337958 247862 338028
rect 247926 337963 247954 338028
rect 247822 337952 247874 337958
rect 247822 337894 247874 337900
rect 247912 337954 247968 337963
rect 247912 337889 247968 337898
rect 248018 337890 248046 338028
rect 248110 337890 248138 338028
rect 248006 337884 248058 337890
rect 248006 337826 248058 337832
rect 248098 337884 248150 337890
rect 248098 337826 248150 337832
rect 247868 337816 247920 337822
rect 247868 337758 247920 337764
rect 247958 337784 248014 337793
rect 247696 337708 247770 337736
rect 247592 337680 247644 337686
rect 247592 337622 247644 337628
rect 247500 336320 247552 336326
rect 247500 336262 247552 336268
rect 247406 333160 247462 333169
rect 247406 333095 247462 333104
rect 247408 333056 247460 333062
rect 247408 332998 247460 333004
rect 247316 320816 247368 320822
rect 247316 320758 247368 320764
rect 247224 10532 247276 10538
rect 247224 10474 247276 10480
rect 247328 10402 247356 320758
rect 247420 11762 247448 332998
rect 247604 331906 247632 337622
rect 247592 331900 247644 331906
rect 247592 331842 247644 331848
rect 247696 328454 247724 337708
rect 247776 337612 247828 337618
rect 247776 337554 247828 337560
rect 247788 336462 247816 337554
rect 247776 336456 247828 336462
rect 247776 336398 247828 336404
rect 247776 333192 247828 333198
rect 247776 333134 247828 333140
rect 247512 328426 247724 328454
rect 247512 153882 247540 328426
rect 247788 316034 247816 333134
rect 247880 332874 247908 337758
rect 248202 337770 248230 338028
rect 248294 337958 248322 338028
rect 248386 337958 248414 338028
rect 248282 337952 248334 337958
rect 248282 337894 248334 337900
rect 248374 337952 248426 337958
rect 248374 337894 248426 337900
rect 248478 337890 248506 338028
rect 248570 337929 248598 338028
rect 248662 337958 248690 338028
rect 248754 337958 248782 338028
rect 248846 337958 248874 338028
rect 248938 337958 248966 338028
rect 248650 337952 248702 337958
rect 248556 337920 248612 337929
rect 248466 337884 248518 337890
rect 248650 337894 248702 337900
rect 248742 337952 248794 337958
rect 248742 337894 248794 337900
rect 248834 337952 248886 337958
rect 248834 337894 248886 337900
rect 248926 337952 248978 337958
rect 248926 337894 248978 337900
rect 248556 337855 248612 337864
rect 248466 337826 248518 337832
rect 248788 337816 248840 337822
rect 247958 337719 248014 337728
rect 248064 337742 248230 337770
rect 248694 337784 248750 337793
rect 248512 337748 248564 337754
rect 247972 333062 248000 337719
rect 248064 333266 248092 337742
rect 248788 337758 248840 337764
rect 248694 337719 248750 337728
rect 248512 337690 248564 337696
rect 248328 337680 248380 337686
rect 248328 337622 248380 337628
rect 248236 337544 248288 337550
rect 248236 337486 248288 337492
rect 248144 337476 248196 337482
rect 248144 337418 248196 337424
rect 248052 333260 248104 333266
rect 248052 333202 248104 333208
rect 247960 333056 248012 333062
rect 247960 332998 248012 333004
rect 247880 332846 248000 332874
rect 247868 330540 247920 330546
rect 247868 330482 247920 330488
rect 247696 316006 247816 316034
rect 247696 160750 247724 316006
rect 247684 160744 247736 160750
rect 247684 160686 247736 160692
rect 247592 159792 247644 159798
rect 247592 159734 247644 159740
rect 247500 153876 247552 153882
rect 247500 153818 247552 153824
rect 247408 11756 247460 11762
rect 247408 11698 247460 11704
rect 247316 10396 247368 10402
rect 247316 10338 247368 10344
rect 246856 6588 246908 6594
rect 246856 6530 246908 6536
rect 246212 4888 246264 4894
rect 246212 4830 246264 4836
rect 244924 3596 244976 3602
rect 244924 3538 244976 3544
rect 243464 3454 244136 3482
rect 244844 3454 245240 3482
rect 244108 480 244136 3454
rect 245212 480 245240 3454
rect 246396 3460 246448 3466
rect 246396 3402 246448 3408
rect 246408 480 246436 3402
rect 247604 480 247632 159734
rect 247880 9353 247908 330482
rect 247866 9344 247922 9353
rect 247866 9279 247922 9288
rect 247972 9217 248000 332846
rect 248156 329186 248184 337418
rect 248144 329180 248196 329186
rect 248144 329122 248196 329128
rect 248248 329118 248276 337486
rect 248340 330546 248368 337622
rect 248420 336660 248472 336666
rect 248420 336602 248472 336608
rect 248432 335850 248460 336602
rect 248420 335844 248472 335850
rect 248420 335786 248472 335792
rect 248524 333305 248552 337690
rect 248604 337680 248656 337686
rect 248604 337622 248656 337628
rect 248616 336394 248644 337622
rect 248604 336388 248656 336394
rect 248604 336330 248656 336336
rect 248708 336274 248736 337719
rect 248616 336246 248736 336274
rect 248510 333296 248566 333305
rect 248510 333231 248566 333240
rect 248328 330540 248380 330546
rect 248328 330482 248380 330488
rect 248236 329112 248288 329118
rect 248236 329054 248288 329060
rect 248326 158264 248382 158273
rect 248326 158199 248382 158208
rect 248234 153776 248290 153785
rect 248234 153711 248290 153720
rect 247958 9208 248014 9217
rect 247958 9143 248014 9152
rect 248248 6526 248276 153711
rect 248340 6730 248368 158199
rect 248616 9489 248644 336246
rect 248800 333198 248828 337758
rect 248880 337748 248932 337754
rect 249030 337736 249058 338028
rect 249122 337958 249150 338028
rect 249214 337958 249242 338028
rect 249306 337958 249334 338028
rect 249110 337952 249162 337958
rect 249110 337894 249162 337900
rect 249202 337952 249254 337958
rect 249202 337894 249254 337900
rect 249294 337952 249346 337958
rect 249294 337894 249346 337900
rect 249398 337770 249426 338028
rect 249490 337822 249518 338028
rect 249582 337963 249610 338028
rect 249568 337954 249624 337963
rect 249674 337958 249702 338028
rect 249766 337958 249794 338028
rect 249858 337958 249886 338028
rect 249568 337889 249624 337898
rect 249662 337952 249714 337958
rect 249662 337894 249714 337900
rect 249754 337952 249806 337958
rect 249754 337894 249806 337900
rect 249846 337952 249898 337958
rect 249950 337929 249978 338028
rect 250042 337958 250070 338028
rect 250134 337958 250162 338028
rect 250226 337958 250254 338028
rect 250030 337952 250082 337958
rect 249846 337894 249898 337900
rect 249936 337920 249992 337929
rect 250030 337894 250082 337900
rect 250122 337952 250174 337958
rect 250122 337894 250174 337900
rect 250214 337952 250266 337958
rect 250214 337894 250266 337900
rect 249936 337855 249992 337864
rect 249352 337742 249426 337770
rect 249478 337816 249530 337822
rect 249478 337758 249530 337764
rect 249984 337816 250036 337822
rect 250214 337816 250266 337822
rect 249984 337758 250036 337764
rect 250212 337784 250214 337793
rect 250266 337784 250268 337793
rect 249616 337748 249668 337754
rect 249030 337708 249104 337736
rect 248880 337690 248932 337696
rect 248892 334778 248920 337690
rect 248972 337340 249024 337346
rect 248972 337282 249024 337288
rect 248984 337074 249012 337282
rect 248972 337068 249024 337074
rect 248972 337010 249024 337016
rect 248972 336252 249024 336258
rect 248972 336194 249024 336200
rect 248984 335850 249012 336194
rect 248972 335844 249024 335850
rect 248972 335786 249024 335792
rect 248972 335708 249024 335714
rect 248972 335650 249024 335656
rect 248984 334966 249012 335650
rect 248972 334960 249024 334966
rect 248972 334902 249024 334908
rect 248892 334750 249012 334778
rect 248880 334552 248932 334558
rect 248880 334494 248932 334500
rect 248788 333192 248840 333198
rect 248788 333134 248840 333140
rect 248696 333124 248748 333130
rect 248696 333066 248748 333072
rect 248708 177410 248736 333066
rect 248788 333056 248840 333062
rect 248788 332998 248840 333004
rect 248800 177478 248828 332998
rect 248892 178770 248920 334494
rect 248984 331809 249012 334750
rect 248970 331800 249026 331809
rect 248970 331735 249026 331744
rect 248972 331696 249024 331702
rect 248972 331638 249024 331644
rect 248880 178764 248932 178770
rect 248880 178706 248932 178712
rect 248788 177472 248840 177478
rect 248788 177414 248840 177420
rect 248696 177404 248748 177410
rect 248696 177346 248748 177352
rect 248696 160540 248748 160546
rect 248696 160482 248748 160488
rect 248708 16574 248736 160482
rect 248708 16546 248828 16574
rect 248602 9480 248658 9489
rect 248602 9415 248658 9424
rect 248328 6724 248380 6730
rect 248328 6666 248380 6672
rect 248236 6520 248288 6526
rect 248236 6462 248288 6468
rect 248800 480 248828 16546
rect 248984 4962 249012 331638
rect 249076 327758 249104 337708
rect 249156 337680 249208 337686
rect 249156 337622 249208 337628
rect 249352 337634 249380 337742
rect 249616 337690 249668 337696
rect 249430 337648 249486 337657
rect 249168 334558 249196 337622
rect 249248 337612 249300 337618
rect 249352 337606 249430 337634
rect 249430 337583 249486 337592
rect 249524 337612 249576 337618
rect 249248 337554 249300 337560
rect 249524 337554 249576 337560
rect 249260 334966 249288 337554
rect 249340 337544 249392 337550
rect 249340 337486 249392 337492
rect 249248 334960 249300 334966
rect 249248 334902 249300 334908
rect 249248 334620 249300 334626
rect 249248 334562 249300 334568
rect 249156 334552 249208 334558
rect 249156 334494 249208 334500
rect 249156 334416 249208 334422
rect 249156 334358 249208 334364
rect 249064 327752 249116 327758
rect 249064 327694 249116 327700
rect 249168 327570 249196 334358
rect 249076 327542 249196 327570
rect 248972 4956 249024 4962
rect 248972 4898 249024 4904
rect 249076 3806 249104 327542
rect 249260 316034 249288 334562
rect 249352 325694 249380 337486
rect 249432 334960 249484 334966
rect 249432 334902 249484 334908
rect 249444 333130 249472 334902
rect 249432 333124 249484 333130
rect 249432 333066 249484 333072
rect 249536 329225 249564 337554
rect 249628 333062 249656 337690
rect 249708 337680 249760 337686
rect 249708 337622 249760 337628
rect 249616 333056 249668 333062
rect 249616 332998 249668 333004
rect 249720 331702 249748 337622
rect 249892 337544 249944 337550
rect 249996 337521 250024 337758
rect 250212 337719 250268 337728
rect 250318 337736 250346 338028
rect 250410 337963 250438 338028
rect 250396 337954 250452 337963
rect 250396 337889 250452 337898
rect 250502 337736 250530 338028
rect 250594 337890 250622 338028
rect 250582 337884 250634 337890
rect 250582 337826 250634 337832
rect 250686 337736 250714 338028
rect 250778 337958 250806 338028
rect 250870 337958 250898 338028
rect 250962 337963 250990 338028
rect 250766 337952 250818 337958
rect 250766 337894 250818 337900
rect 250858 337952 250910 337958
rect 250858 337894 250910 337900
rect 250948 337954 251004 337963
rect 251054 337958 251082 338028
rect 250948 337889 251004 337898
rect 251042 337952 251094 337958
rect 251042 337894 251094 337900
rect 251146 337890 251174 338028
rect 251238 337963 251266 338028
rect 251224 337954 251280 337963
rect 251134 337884 251186 337890
rect 251224 337889 251280 337898
rect 251330 337890 251358 338028
rect 251422 337958 251450 338028
rect 251410 337952 251462 337958
rect 251410 337894 251462 337900
rect 251134 337826 251186 337832
rect 251318 337884 251370 337890
rect 251318 337826 251370 337832
rect 250318 337708 250392 337736
rect 250258 337648 250314 337657
rect 250258 337583 250314 337592
rect 249892 337486 249944 337492
rect 249982 337512 250038 337521
rect 249800 336932 249852 336938
rect 249800 336874 249852 336880
rect 249812 336394 249840 336874
rect 249800 336388 249852 336394
rect 249800 336330 249852 336336
rect 249708 331696 249760 331702
rect 249708 331638 249760 331644
rect 249522 329216 249578 329225
rect 249522 329151 249578 329160
rect 249352 325666 249564 325694
rect 249168 316006 249288 316034
rect 249168 6322 249196 316006
rect 249536 7614 249564 325666
rect 249708 158636 249760 158642
rect 249708 158578 249760 158584
rect 249616 158500 249668 158506
rect 249616 158442 249668 158448
rect 249524 7608 249576 7614
rect 249524 7550 249576 7556
rect 249628 6322 249656 158442
rect 249156 6316 249208 6322
rect 249156 6258 249208 6264
rect 249616 6316 249668 6322
rect 249616 6258 249668 6264
rect 249720 4078 249748 158578
rect 249904 6225 249932 337486
rect 249982 337447 250038 337456
rect 250168 337068 250220 337074
rect 250168 337010 250220 337016
rect 250076 333260 250128 333266
rect 250076 333202 250128 333208
rect 249984 333192 250036 333198
rect 249984 333134 250036 333140
rect 249996 6254 250024 333134
rect 250088 9586 250116 333202
rect 250180 10470 250208 337010
rect 250272 333266 250300 337583
rect 250364 337482 250392 337708
rect 250456 337708 250530 337736
rect 250640 337708 250714 337736
rect 251180 337748 251232 337754
rect 250352 337476 250404 337482
rect 250352 337418 250404 337424
rect 250260 333260 250312 333266
rect 250260 333202 250312 333208
rect 250352 333260 250404 333266
rect 250352 333202 250404 333208
rect 250260 333124 250312 333130
rect 250260 333066 250312 333072
rect 250272 11830 250300 333066
rect 250364 12306 250392 333202
rect 250456 177546 250484 337708
rect 250536 337612 250588 337618
rect 250536 337554 250588 337560
rect 250548 178838 250576 337554
rect 250640 337074 250668 337708
rect 251514 337736 251542 338028
rect 251606 337929 251634 338028
rect 251698 337958 251726 338028
rect 251686 337952 251738 337958
rect 251592 337920 251648 337929
rect 251686 337894 251738 337900
rect 251592 337855 251648 337864
rect 251640 337816 251692 337822
rect 251640 337758 251692 337764
rect 251790 337770 251818 338028
rect 251882 337890 251910 338028
rect 251974 337963 252002 338028
rect 251960 337954 252016 337963
rect 252066 337958 252094 338028
rect 251870 337884 251922 337890
rect 251960 337889 252016 337898
rect 252054 337952 252106 337958
rect 252054 337894 252106 337900
rect 251870 337826 251922 337832
rect 252008 337816 252060 337822
rect 251914 337784 251970 337793
rect 251180 337690 251232 337696
rect 251284 337708 251542 337736
rect 250996 337680 251048 337686
rect 250996 337622 251048 337628
rect 250720 337612 250772 337618
rect 250720 337554 250772 337560
rect 250628 337068 250680 337074
rect 250628 337010 250680 337016
rect 250732 333266 250760 337554
rect 250810 337512 250866 337521
rect 250810 337447 250866 337456
rect 250904 337476 250956 337482
rect 250720 333260 250772 333266
rect 250720 333202 250772 333208
rect 250824 333198 250852 337447
rect 250904 337418 250956 337424
rect 250812 333192 250864 333198
rect 250812 333134 250864 333140
rect 250916 316034 250944 337418
rect 251008 333130 251036 337622
rect 251088 337612 251140 337618
rect 251088 337554 251140 337560
rect 251100 337385 251128 337554
rect 251086 337376 251142 337385
rect 251086 337311 251142 337320
rect 250996 333124 251048 333130
rect 250996 333066 251048 333072
rect 251192 331974 251220 337690
rect 251284 333305 251312 337708
rect 251364 337612 251416 337618
rect 251364 337554 251416 337560
rect 251548 337612 251600 337618
rect 251548 337554 251600 337560
rect 251376 334626 251404 337554
rect 251456 337544 251508 337550
rect 251456 337486 251508 337492
rect 251364 334620 251416 334626
rect 251364 334562 251416 334568
rect 251468 333441 251496 337486
rect 251454 333432 251510 333441
rect 251454 333367 251510 333376
rect 251560 333334 251588 337554
rect 251652 337278 251680 337758
rect 251790 337742 251864 337770
rect 251732 337612 251784 337618
rect 251732 337554 251784 337560
rect 251640 337272 251692 337278
rect 251640 337214 251692 337220
rect 251548 333328 251600 333334
rect 251270 333296 251326 333305
rect 251548 333270 251600 333276
rect 251270 333231 251326 333240
rect 251180 331968 251232 331974
rect 251180 331910 251232 331916
rect 251640 331016 251692 331022
rect 251640 330958 251692 330964
rect 251180 330948 251232 330954
rect 251180 330890 251232 330896
rect 251192 330682 251220 330890
rect 251180 330676 251232 330682
rect 251180 330618 251232 330624
rect 251364 330676 251416 330682
rect 251364 330618 251416 330624
rect 250824 316006 250944 316034
rect 250536 178832 250588 178838
rect 250536 178774 250588 178780
rect 250444 177540 250496 177546
rect 250444 177482 250496 177488
rect 250444 156936 250496 156942
rect 250444 156878 250496 156884
rect 250352 12300 250404 12306
rect 250352 12242 250404 12248
rect 250260 11824 250312 11830
rect 250260 11766 250312 11772
rect 250168 10464 250220 10470
rect 250168 10406 250220 10412
rect 250076 9580 250128 9586
rect 250076 9522 250128 9528
rect 249984 6248 250036 6254
rect 249890 6216 249946 6225
rect 249984 6190 250036 6196
rect 249890 6151 249946 6160
rect 249708 4072 249760 4078
rect 249708 4014 249760 4020
rect 249064 3800 249116 3806
rect 249064 3742 249116 3748
rect 240478 354 240590 480
rect 240152 326 240590 354
rect 240478 -960 240590 326
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 354 250066 480
rect 250456 354 250484 156878
rect 250824 5030 250852 316006
rect 250996 160744 251048 160750
rect 250996 160686 251048 160692
rect 251008 6254 251036 160686
rect 251088 158568 251140 158574
rect 251088 158510 251140 158516
rect 250996 6248 251048 6254
rect 250996 6190 251048 6196
rect 250812 5024 250864 5030
rect 250812 4966 250864 4972
rect 251100 3942 251128 158510
rect 251376 10742 251404 330618
rect 251548 330540 251600 330546
rect 251548 330482 251600 330488
rect 251456 330472 251508 330478
rect 251456 330414 251508 330420
rect 251468 11966 251496 330414
rect 251560 82142 251588 330482
rect 251652 330342 251680 330958
rect 251640 330336 251692 330342
rect 251640 330278 251692 330284
rect 251640 159860 251692 159866
rect 251640 159802 251692 159808
rect 251548 82136 251600 82142
rect 251548 82078 251600 82084
rect 251456 11960 251508 11966
rect 251456 11902 251508 11908
rect 251364 10736 251416 10742
rect 251364 10678 251416 10684
rect 251652 6914 251680 159802
rect 251192 6886 251680 6914
rect 251088 3936 251140 3942
rect 251088 3878 251140 3884
rect 251192 480 251220 6886
rect 251744 6361 251772 337554
rect 251836 330562 251864 337742
rect 252008 337758 252060 337764
rect 252158 337770 252186 338028
rect 252250 337890 252278 338028
rect 252342 337958 252370 338028
rect 252434 337963 252462 338028
rect 252330 337952 252382 337958
rect 252330 337894 252382 337900
rect 252420 337954 252476 337963
rect 252238 337884 252290 337890
rect 252420 337889 252476 337898
rect 252238 337826 252290 337832
rect 252282 337784 252338 337793
rect 251914 337719 251970 337728
rect 251928 335918 251956 337719
rect 251916 335912 251968 335918
rect 251916 335854 251968 335860
rect 251916 335640 251968 335646
rect 251916 335582 251968 335588
rect 251928 331022 251956 335582
rect 251916 331016 251968 331022
rect 251916 330958 251968 330964
rect 252020 330682 252048 337758
rect 252158 337742 252232 337770
rect 252204 335560 252232 337742
rect 252526 337736 252554 338028
rect 252618 337890 252646 338028
rect 252606 337884 252658 337890
rect 252606 337826 252658 337832
rect 252710 337770 252738 338028
rect 252802 337793 252830 338028
rect 252894 337929 252922 338028
rect 252880 337920 252936 337929
rect 252880 337855 252936 337864
rect 252282 337719 252338 337728
rect 252112 335532 252232 335560
rect 252008 330676 252060 330682
rect 252008 330618 252060 330624
rect 251836 330534 252048 330562
rect 252112 330546 252140 335532
rect 252192 335436 252244 335442
rect 252192 335378 252244 335384
rect 251824 330336 251876 330342
rect 251824 330278 251876 330284
rect 251836 9110 251864 330278
rect 252020 325694 252048 330534
rect 252100 330540 252152 330546
rect 252100 330482 252152 330488
rect 252204 327826 252232 335378
rect 252296 333402 252324 337719
rect 252480 337708 252554 337736
rect 252664 337742 252738 337770
rect 252788 337784 252844 337793
rect 252376 337680 252428 337686
rect 252376 337622 252428 337628
rect 252284 333396 252336 333402
rect 252284 333338 252336 333344
rect 252388 330478 252416 337622
rect 252480 335782 252508 337708
rect 252560 337612 252612 337618
rect 252560 337554 252612 337560
rect 252468 335776 252520 335782
rect 252468 335718 252520 335724
rect 252468 335572 252520 335578
rect 252468 335514 252520 335520
rect 252480 330954 252508 335514
rect 252468 330948 252520 330954
rect 252468 330890 252520 330896
rect 252572 330546 252600 337554
rect 252664 334801 252692 337742
rect 252986 337770 253014 338028
rect 253078 337929 253106 338028
rect 253064 337920 253120 337929
rect 253170 337890 253198 338028
rect 253262 337890 253290 338028
rect 253064 337855 253120 337864
rect 253158 337884 253210 337890
rect 253158 337826 253210 337832
rect 253250 337884 253302 337890
rect 253250 337826 253302 337832
rect 253202 337784 253258 337793
rect 252986 337742 253060 337770
rect 252788 337719 252844 337728
rect 252836 337612 252888 337618
rect 252836 337554 252888 337560
rect 252650 334792 252706 334801
rect 252650 334727 252706 334736
rect 252848 331214 252876 337554
rect 252756 331186 252876 331214
rect 252560 330540 252612 330546
rect 252560 330482 252612 330488
rect 252376 330472 252428 330478
rect 252376 330414 252428 330420
rect 252652 330404 252704 330410
rect 252652 330346 252704 330352
rect 252192 327820 252244 327826
rect 252192 327762 252244 327768
rect 252020 325666 252140 325694
rect 251824 9104 251876 9110
rect 251824 9046 251876 9052
rect 252112 7682 252140 325666
rect 252664 12170 252692 330346
rect 252652 12164 252704 12170
rect 252652 12106 252704 12112
rect 252756 12034 252784 331186
rect 253032 330970 253060 337742
rect 253354 337770 253382 338028
rect 253446 337958 253474 338028
rect 253434 337952 253486 337958
rect 253434 337894 253486 337900
rect 253538 337770 253566 338028
rect 253630 337890 253658 338028
rect 253618 337884 253670 337890
rect 253618 337826 253670 337832
rect 253722 337770 253750 338028
rect 253354 337742 253428 337770
rect 253202 337719 253258 337728
rect 253112 337680 253164 337686
rect 253112 337622 253164 337628
rect 252848 330942 253060 330970
rect 252848 330682 252876 330942
rect 253124 330834 253152 337622
rect 253216 336705 253244 337719
rect 253296 337680 253348 337686
rect 253296 337622 253348 337628
rect 253202 336696 253258 336705
rect 253202 336631 253258 336640
rect 253308 335986 253336 337622
rect 253296 335980 253348 335986
rect 253296 335922 253348 335928
rect 253204 334620 253256 334626
rect 253204 334562 253256 334568
rect 252940 330806 253152 330834
rect 252836 330676 252888 330682
rect 252836 330618 252888 330624
rect 252836 330540 252888 330546
rect 252836 330482 252888 330488
rect 252848 12102 252876 330482
rect 252940 14482 252968 330806
rect 253112 330676 253164 330682
rect 253112 330618 253164 330624
rect 253020 330472 253072 330478
rect 253020 330414 253072 330420
rect 253032 14550 253060 330414
rect 253124 178906 253152 330618
rect 253216 178974 253244 334562
rect 253296 330540 253348 330546
rect 253296 330482 253348 330488
rect 253308 179042 253336 330482
rect 253400 325694 253428 337742
rect 253492 337742 253566 337770
rect 253676 337742 253750 337770
rect 253492 334626 253520 337742
rect 253572 336252 253624 336258
rect 253572 336194 253624 336200
rect 253480 334620 253532 334626
rect 253480 334562 253532 334568
rect 253584 331214 253612 336194
rect 253492 331186 253612 331214
rect 253492 329390 253520 331186
rect 253676 330410 253704 337742
rect 253814 337634 253842 338028
rect 253906 337958 253934 338028
rect 253998 337963 254026 338028
rect 253894 337952 253946 337958
rect 253894 337894 253946 337900
rect 253984 337954 254040 337963
rect 253984 337889 254040 337898
rect 254090 337822 254118 338028
rect 254182 337963 254210 338028
rect 254168 337954 254224 337963
rect 254168 337889 254224 337898
rect 254274 337890 254302 338028
rect 254366 337963 254394 338028
rect 254352 337954 254408 337963
rect 254262 337884 254314 337890
rect 254352 337889 254408 337898
rect 254458 337890 254486 338028
rect 254262 337826 254314 337832
rect 254446 337884 254498 337890
rect 254446 337826 254498 337832
rect 254550 337822 254578 338028
rect 254642 337822 254670 338028
rect 254734 337822 254762 338028
rect 254078 337816 254130 337822
rect 254078 337758 254130 337764
rect 254538 337816 254590 337822
rect 254538 337758 254590 337764
rect 254630 337816 254682 337822
rect 254630 337758 254682 337764
rect 254722 337816 254774 337822
rect 254826 337804 254854 338028
rect 254918 337958 254946 338028
rect 255010 337963 255038 338028
rect 254906 337952 254958 337958
rect 254906 337894 254958 337900
rect 254996 337954 255052 337963
rect 255102 337958 255130 338028
rect 255194 337958 255222 338028
rect 255286 337958 255314 338028
rect 255378 337958 255406 338028
rect 255470 337963 255498 338028
rect 254996 337889 255052 337898
rect 255090 337952 255142 337958
rect 255090 337894 255142 337900
rect 255182 337952 255234 337958
rect 255182 337894 255234 337900
rect 255274 337952 255326 337958
rect 255274 337894 255326 337900
rect 255366 337952 255418 337958
rect 255366 337894 255418 337900
rect 255456 337954 255512 337963
rect 255456 337889 255512 337898
rect 255562 337827 255590 338028
rect 255654 337963 255682 338028
rect 255640 337954 255696 337963
rect 255640 337889 255696 337898
rect 255044 337816 255096 337822
rect 254826 337776 254900 337804
rect 254722 337758 254774 337764
rect 253940 337748 253992 337754
rect 253940 337690 253992 337696
rect 254216 337748 254268 337754
rect 254216 337690 254268 337696
rect 253768 337606 253842 337634
rect 253768 330546 253796 337606
rect 253952 337498 253980 337690
rect 254124 337680 254176 337686
rect 254124 337622 254176 337628
rect 253860 337470 253980 337498
rect 253756 330540 253808 330546
rect 253756 330482 253808 330488
rect 253860 330478 253888 337470
rect 253938 337376 253994 337385
rect 253938 337311 253940 337320
rect 253992 337311 253994 337320
rect 253940 337282 253992 337288
rect 253940 334620 253992 334626
rect 253940 334562 253992 334568
rect 253848 330472 253900 330478
rect 253848 330414 253900 330420
rect 253664 330404 253716 330410
rect 253664 330346 253716 330352
rect 253480 329384 253532 329390
rect 253480 329326 253532 329332
rect 253952 329254 253980 334562
rect 254136 334529 254164 337622
rect 254122 334520 254178 334529
rect 254122 334455 254178 334464
rect 254228 332897 254256 337690
rect 254768 337680 254820 337686
rect 254768 337622 254820 337628
rect 254308 337612 254360 337618
rect 254308 337554 254360 337560
rect 254676 337612 254728 337618
rect 254676 337554 254728 337560
rect 254214 332888 254270 332897
rect 254214 332823 254270 332832
rect 254320 331214 254348 337554
rect 254492 337544 254544 337550
rect 254398 337512 254454 337521
rect 254544 337504 254624 337532
rect 254492 337486 254544 337492
rect 254398 337447 254454 337456
rect 254136 331186 254348 331214
rect 253940 329248 253992 329254
rect 253940 329190 253992 329196
rect 253400 325666 253704 325694
rect 253296 179036 253348 179042
rect 253296 178978 253348 178984
rect 253204 178968 253256 178974
rect 253204 178910 253256 178916
rect 253112 178900 253164 178906
rect 253112 178842 253164 178848
rect 253110 158672 253166 158681
rect 253110 158607 253166 158616
rect 253124 16574 253152 158607
rect 253124 16546 253520 16574
rect 253020 14544 253072 14550
rect 253020 14486 253072 14492
rect 252928 14476 252980 14482
rect 252928 14418 252980 14424
rect 252836 12096 252888 12102
rect 252836 12038 252888 12044
rect 252744 12028 252796 12034
rect 252744 11970 252796 11976
rect 252100 7676 252152 7682
rect 252100 7618 252152 7624
rect 251730 6352 251786 6361
rect 251730 6287 251786 6296
rect 252376 3188 252428 3194
rect 252376 3130 252428 3136
rect 252388 480 252416 3130
rect 253492 480 253520 16546
rect 253676 7954 253704 325666
rect 253848 157956 253900 157962
rect 253848 157898 253900 157904
rect 253756 155508 253808 155514
rect 253756 155450 253808 155456
rect 253664 7948 253716 7954
rect 253664 7890 253716 7896
rect 253768 3330 253796 155450
rect 253860 4146 253888 157898
rect 254136 12238 254164 331186
rect 254308 326460 254360 326466
rect 254308 326402 254360 326408
rect 254216 326324 254268 326330
rect 254216 326266 254268 326272
rect 254228 13190 254256 326266
rect 254320 14618 254348 326402
rect 254412 179110 254440 337447
rect 254492 335368 254544 335374
rect 254492 335310 254544 335316
rect 254504 331214 254532 335310
rect 254596 333470 254624 337504
rect 254584 333464 254636 333470
rect 254584 333406 254636 333412
rect 254504 331186 254624 331214
rect 254492 326392 254544 326398
rect 254492 326334 254544 326340
rect 254400 179104 254452 179110
rect 254400 179046 254452 179052
rect 254308 14612 254360 14618
rect 254308 14554 254360 14560
rect 254216 13184 254268 13190
rect 254216 13126 254268 13132
rect 254124 12232 254176 12238
rect 254124 12174 254176 12180
rect 254504 6905 254532 326334
rect 254596 7818 254624 331186
rect 254688 326346 254716 337554
rect 254780 326466 254808 337622
rect 254768 326460 254820 326466
rect 254768 326402 254820 326408
rect 254688 326318 254808 326346
rect 254872 326330 254900 337776
rect 255044 337758 255096 337764
rect 255136 337816 255188 337822
rect 255136 337758 255188 337764
rect 255548 337818 255604 337827
rect 255056 336054 255084 337758
rect 255044 336048 255096 336054
rect 255044 335990 255096 335996
rect 255148 334626 255176 337758
rect 255228 337748 255280 337754
rect 255548 337753 255604 337762
rect 255228 337690 255280 337696
rect 255136 334620 255188 334626
rect 255136 334562 255188 334568
rect 254952 330336 255004 330342
rect 254952 330278 255004 330284
rect 254676 325984 254728 325990
rect 254676 325926 254728 325932
rect 254584 7812 254636 7818
rect 254584 7754 254636 7760
rect 254688 6914 254716 325926
rect 254490 6896 254546 6905
rect 254490 6831 254546 6840
rect 254596 6886 254716 6914
rect 253848 4140 253900 4146
rect 253848 4082 253900 4088
rect 254596 3466 254624 6886
rect 254780 6497 254808 326318
rect 254860 326324 254912 326330
rect 254860 326266 254912 326272
rect 254964 325990 254992 330278
rect 255240 326398 255268 337690
rect 255504 337680 255556 337686
rect 255424 337640 255504 337668
rect 255320 337612 255372 337618
rect 255320 337554 255372 337560
rect 255332 336122 255360 337554
rect 255320 336116 255372 336122
rect 255320 336058 255372 336064
rect 255320 335980 255372 335986
rect 255320 335922 255372 335928
rect 255332 333606 255360 335922
rect 255320 333600 255372 333606
rect 255320 333542 255372 333548
rect 255424 332042 255452 337640
rect 255746 337668 255774 338028
rect 255838 337929 255866 338028
rect 255824 337920 255880 337929
rect 255824 337855 255880 337864
rect 255930 337668 255958 338028
rect 256022 337736 256050 338028
rect 256114 337929 256142 338028
rect 256206 337958 256234 338028
rect 256194 337952 256246 337958
rect 256100 337920 256156 337929
rect 256194 337894 256246 337900
rect 256100 337855 256156 337864
rect 256298 337804 256326 338028
rect 256160 337776 256326 337804
rect 256022 337708 256096 337736
rect 255504 337622 255556 337628
rect 255594 337648 255650 337657
rect 255746 337640 255820 337668
rect 255930 337640 256004 337668
rect 255594 337583 255650 337592
rect 255504 336320 255556 336326
rect 255504 336262 255556 336268
rect 255412 332036 255464 332042
rect 255412 331978 255464 331984
rect 255228 326392 255280 326398
rect 255228 326334 255280 326340
rect 254952 325984 255004 325990
rect 254952 325926 255004 325932
rect 255228 158704 255280 158710
rect 255228 158646 255280 158652
rect 254766 6488 254822 6497
rect 254766 6423 254822 6432
rect 254676 3528 254728 3534
rect 254676 3470 254728 3476
rect 254584 3460 254636 3466
rect 254584 3402 254636 3408
rect 253756 3324 253808 3330
rect 253756 3266 253808 3272
rect 254688 480 254716 3470
rect 255240 3369 255268 158646
rect 255516 8022 255544 336262
rect 255608 333538 255636 337583
rect 255688 337476 255740 337482
rect 255688 337418 255740 337424
rect 255700 335424 255728 337418
rect 255792 335782 255820 337640
rect 255870 337512 255926 337521
rect 255870 337447 255926 337456
rect 255780 335776 255832 335782
rect 255780 335718 255832 335724
rect 255884 335646 255912 337447
rect 255976 335889 256004 337640
rect 255962 335880 256018 335889
rect 255962 335815 256018 335824
rect 255964 335776 256016 335782
rect 255964 335718 256016 335724
rect 255872 335640 255924 335646
rect 255872 335582 255924 335588
rect 255700 335396 255820 335424
rect 255688 335300 255740 335306
rect 255688 335242 255740 335248
rect 255596 333532 255648 333538
rect 255596 333474 255648 333480
rect 255700 332594 255728 335242
rect 255608 332566 255728 332594
rect 255608 21418 255636 332566
rect 255792 326346 255820 335396
rect 255976 334762 256004 335718
rect 256068 334830 256096 337708
rect 256056 334824 256108 334830
rect 256056 334766 256108 334772
rect 255964 334756 256016 334762
rect 255964 334698 256016 334704
rect 256160 331214 256188 337776
rect 256390 337668 256418 338028
rect 256482 337736 256510 338028
rect 256574 337895 256602 338028
rect 256560 337886 256616 337895
rect 256666 337890 256694 338028
rect 256758 337963 256786 338028
rect 256744 337954 256800 337963
rect 256560 337821 256616 337830
rect 256654 337884 256706 337890
rect 256744 337889 256800 337898
rect 256850 337890 256878 338028
rect 256654 337826 256706 337832
rect 256838 337884 256890 337890
rect 256838 337826 256890 337832
rect 256942 337736 256970 338028
rect 256482 337708 256648 337736
rect 256344 337640 256418 337668
rect 256514 337648 256570 337657
rect 256344 335306 256372 337640
rect 256514 337583 256570 337592
rect 256424 337544 256476 337550
rect 256424 337486 256476 337492
rect 256436 336734 256464 337486
rect 256424 336728 256476 336734
rect 256424 336670 256476 336676
rect 256424 336048 256476 336054
rect 256424 335990 256476 335996
rect 256332 335300 256384 335306
rect 256332 335242 256384 335248
rect 256436 333690 256464 335990
rect 256344 333662 256464 333690
rect 256240 333396 256292 333402
rect 256240 333338 256292 333344
rect 255700 326318 255820 326346
rect 255884 331186 256188 331214
rect 255700 177614 255728 326318
rect 255884 321554 255912 331186
rect 255964 330676 256016 330682
rect 255964 330618 256016 330624
rect 255792 321526 255912 321554
rect 255688 177608 255740 177614
rect 255688 177550 255740 177556
rect 255686 159488 255742 159497
rect 255686 159423 255742 159432
rect 255596 21412 255648 21418
rect 255596 21354 255648 21360
rect 255504 8016 255556 8022
rect 255504 7958 255556 7964
rect 255700 3482 255728 159423
rect 255792 5166 255820 321526
rect 255780 5160 255832 5166
rect 255780 5102 255832 5108
rect 255700 3454 255912 3482
rect 255226 3360 255282 3369
rect 255226 3295 255282 3304
rect 255884 480 255912 3454
rect 255976 3194 256004 330618
rect 256148 326460 256200 326466
rect 256148 326402 256200 326408
rect 256054 326360 256110 326369
rect 256054 326295 256110 326304
rect 256068 3534 256096 326295
rect 256160 6633 256188 326402
rect 256252 326074 256280 333338
rect 256344 326262 256372 333662
rect 256424 333600 256476 333606
rect 256424 333542 256476 333548
rect 256436 326346 256464 333542
rect 256528 326466 256556 337583
rect 256620 336326 256648 337708
rect 256712 337708 256970 337736
rect 256608 336320 256660 336326
rect 256608 336262 256660 336268
rect 256712 333878 256740 337708
rect 256792 337612 256844 337618
rect 257034 337600 257062 338028
rect 257126 337736 257154 338028
rect 257218 337804 257246 338028
rect 257310 337958 257338 338028
rect 257402 337958 257430 338028
rect 257298 337952 257350 337958
rect 257298 337894 257350 337900
rect 257390 337952 257442 337958
rect 257494 337929 257522 338028
rect 257586 337958 257614 338028
rect 257574 337952 257626 337958
rect 257390 337894 257442 337900
rect 257480 337920 257536 337929
rect 257574 337894 257626 337900
rect 257678 337890 257706 338028
rect 257770 337929 257798 338028
rect 257756 337920 257812 337929
rect 257480 337855 257536 337864
rect 257666 337884 257718 337890
rect 257756 337855 257812 337864
rect 257666 337826 257718 337832
rect 257862 337822 257890 338028
rect 257954 337958 257982 338028
rect 257942 337952 257994 337958
rect 257942 337894 257994 337900
rect 257850 337816 257902 337822
rect 257218 337776 257292 337804
rect 257126 337708 257200 337736
rect 257034 337572 257108 337600
rect 256792 337554 256844 337560
rect 256804 334665 256832 337554
rect 256976 337476 257028 337482
rect 256976 337418 257028 337424
rect 256884 337408 256936 337414
rect 256884 337350 256936 337356
rect 256790 334656 256846 334665
rect 256790 334591 256846 334600
rect 256700 333872 256752 333878
rect 256700 333814 256752 333820
rect 256516 326460 256568 326466
rect 256516 326402 256568 326408
rect 256436 326318 256648 326346
rect 256332 326256 256384 326262
rect 256332 326198 256384 326204
rect 256252 326046 256556 326074
rect 256424 325984 256476 325990
rect 256424 325926 256476 325932
rect 256436 163742 256464 325926
rect 256424 163736 256476 163742
rect 256424 163678 256476 163684
rect 256528 100094 256556 326046
rect 256516 100088 256568 100094
rect 256516 100030 256568 100036
rect 256146 6624 256202 6633
rect 256146 6559 256202 6568
rect 256620 3602 256648 326318
rect 256896 177750 256924 337350
rect 256988 329322 257016 337418
rect 257080 335345 257108 337572
rect 257066 335336 257122 335345
rect 257066 335271 257122 335280
rect 257172 334898 257200 337708
rect 257160 334892 257212 334898
rect 257160 334834 257212 334840
rect 257264 331226 257292 337776
rect 257618 337784 257674 337793
rect 257436 337748 257488 337754
rect 258046 337804 258074 338028
rect 258138 337822 258166 338028
rect 257850 337758 257902 337764
rect 258000 337776 258074 337804
rect 258126 337816 258178 337822
rect 257618 337719 257674 337728
rect 257436 337690 257488 337696
rect 257344 337612 257396 337618
rect 257344 337554 257396 337560
rect 257356 334801 257384 337554
rect 257342 334792 257398 334801
rect 257342 334727 257398 334736
rect 257448 334642 257476 337690
rect 257526 337648 257582 337657
rect 257526 337583 257582 337592
rect 257356 334614 257476 334642
rect 257252 331220 257304 331226
rect 257252 331162 257304 331168
rect 256976 329316 257028 329322
rect 256976 329258 257028 329264
rect 257356 327026 257384 334614
rect 257540 333674 257568 337583
rect 257632 334642 257660 337719
rect 257804 337680 257856 337686
rect 257804 337622 257856 337628
rect 257816 336190 257844 337622
rect 257896 337612 257948 337618
rect 257896 337554 257948 337560
rect 257908 337006 257936 337554
rect 257896 337000 257948 337006
rect 257896 336942 257948 336948
rect 257804 336184 257856 336190
rect 257804 336126 257856 336132
rect 257896 336184 257948 336190
rect 257896 336126 257948 336132
rect 257908 335238 257936 336126
rect 257896 335232 257948 335238
rect 257896 335174 257948 335180
rect 257632 334614 257752 334642
rect 257618 333976 257674 333985
rect 257618 333911 257674 333920
rect 257528 333668 257580 333674
rect 257528 333610 257580 333616
rect 257436 333600 257488 333606
rect 257436 333542 257488 333548
rect 257080 326998 257384 327026
rect 256976 326392 257028 326398
rect 256976 326334 257028 326340
rect 256988 179178 257016 326334
rect 257080 191146 257108 326998
rect 257160 326732 257212 326738
rect 257160 326674 257212 326680
rect 257068 191140 257120 191146
rect 257068 191082 257120 191088
rect 256976 179172 257028 179178
rect 256976 179114 257028 179120
rect 257172 177818 257200 326674
rect 257448 326618 257476 333542
rect 257528 331220 257580 331226
rect 257528 331162 257580 331168
rect 257356 326590 257476 326618
rect 257356 321554 257384 326590
rect 257264 321526 257384 321554
rect 257160 177812 257212 177818
rect 257160 177754 257212 177760
rect 256884 177744 256936 177750
rect 256884 177686 256936 177692
rect 256792 157820 256844 157826
rect 256792 157762 256844 157768
rect 256700 153196 256752 153202
rect 256700 153138 256752 153144
rect 256712 152425 256740 153138
rect 256698 152416 256754 152425
rect 256698 152351 256754 152360
rect 256700 144900 256752 144906
rect 256700 144842 256752 144848
rect 256712 143585 256740 144842
rect 256698 143576 256754 143585
rect 256698 143511 256754 143520
rect 256804 142154 256832 157762
rect 257264 148345 257292 321526
rect 257540 316034 257568 331162
rect 257632 326602 257660 333911
rect 257620 326596 257672 326602
rect 257620 326538 257672 326544
rect 257724 326398 257752 334614
rect 257894 332208 257950 332217
rect 257804 332172 257856 332178
rect 257894 332143 257950 332152
rect 257804 332114 257856 332120
rect 257712 326392 257764 326398
rect 257712 326334 257764 326340
rect 257448 316006 257568 316034
rect 257448 177682 257476 316006
rect 257436 177676 257488 177682
rect 257436 177618 257488 177624
rect 257342 163432 257398 163441
rect 257342 163367 257398 163376
rect 257250 148336 257306 148345
rect 257250 148271 257306 148280
rect 256712 142126 256832 142154
rect 256608 3596 256660 3602
rect 256608 3538 256660 3544
rect 256056 3528 256108 3534
rect 256056 3470 256108 3476
rect 255964 3188 256016 3194
rect 255964 3130 256016 3136
rect 249954 326 250484 354
rect 249954 -960 250066 326
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 256712 354 256740 142126
rect 257252 142112 257304 142118
rect 257252 142054 257304 142060
rect 257264 139505 257292 142054
rect 257250 139496 257306 139505
rect 257250 139431 257306 139440
rect 256792 135244 256844 135250
rect 256792 135186 256844 135192
rect 256804 134745 256832 135186
rect 256790 134736 256846 134745
rect 256790 134671 256846 134680
rect 256792 131096 256844 131102
rect 256792 131038 256844 131044
rect 256804 130665 256832 131038
rect 256790 130656 256846 130665
rect 256790 130591 256846 130600
rect 256792 126948 256844 126954
rect 256792 126890 256844 126896
rect 256804 125905 256832 126890
rect 256790 125896 256846 125905
rect 256790 125831 256846 125840
rect 256792 122800 256844 122806
rect 256792 122742 256844 122748
rect 256804 121825 256832 122742
rect 256790 121816 256846 121825
rect 256790 121751 256846 121760
rect 256792 113144 256844 113150
rect 256792 113086 256844 113092
rect 256804 112985 256832 113086
rect 256790 112976 256846 112985
rect 256790 112911 256846 112920
rect 256792 104848 256844 104854
rect 256792 104790 256844 104796
rect 256804 104145 256832 104790
rect 256790 104136 256846 104145
rect 256790 104071 256846 104080
rect 257356 97646 257384 163367
rect 257434 155952 257490 155961
rect 257434 155887 257490 155896
rect 257344 97640 257396 97646
rect 257344 97582 257396 97588
rect 257448 3466 257476 155887
rect 257712 155644 257764 155650
rect 257712 155586 257764 155592
rect 257528 155576 257580 155582
rect 257528 155518 257580 155524
rect 257540 3534 257568 155518
rect 257618 155136 257674 155145
rect 257618 155071 257674 155080
rect 257632 3874 257660 155071
rect 257620 3868 257672 3874
rect 257620 3810 257672 3816
rect 257724 3806 257752 155586
rect 257816 142118 257844 332114
rect 257804 142112 257856 142118
rect 257804 142054 257856 142060
rect 257802 141944 257858 141953
rect 257802 141879 257858 141888
rect 257816 132569 257844 141879
rect 257802 132560 257858 132569
rect 257802 132495 257858 132504
rect 257802 132424 257858 132433
rect 257802 132359 257858 132368
rect 257816 122913 257844 132359
rect 257802 122904 257858 122913
rect 257802 122839 257858 122848
rect 257802 122768 257858 122777
rect 257802 122703 257858 122712
rect 257816 113257 257844 122703
rect 257802 113248 257858 113257
rect 257802 113183 257858 113192
rect 257802 113112 257858 113121
rect 257802 113047 257858 113056
rect 257816 103601 257844 113047
rect 257802 103592 257858 103601
rect 257802 103527 257858 103536
rect 257802 103456 257858 103465
rect 257802 103391 257858 103400
rect 257816 93945 257844 103391
rect 257908 97782 257936 332143
rect 258000 326738 258028 337776
rect 258230 337793 258258 338028
rect 258322 337929 258350 338028
rect 258414 337958 258442 338028
rect 258506 337958 258534 338028
rect 258402 337952 258454 337958
rect 258308 337920 258364 337929
rect 258402 337894 258454 337900
rect 258494 337952 258546 337958
rect 258494 337894 258546 337900
rect 258308 337855 258364 337864
rect 258448 337816 258500 337822
rect 258126 337758 258178 337764
rect 258216 337784 258272 337793
rect 258448 337758 258500 337764
rect 258216 337719 258272 337728
rect 258080 337680 258132 337686
rect 258080 337622 258132 337628
rect 258356 337680 258408 337686
rect 258356 337622 258408 337628
rect 258092 336025 258120 337622
rect 258264 337544 258316 337550
rect 258264 337486 258316 337492
rect 258276 336161 258304 337486
rect 258368 336569 258396 337622
rect 258354 336560 258410 336569
rect 258354 336495 258410 336504
rect 258460 336410 258488 337758
rect 258598 337736 258626 338028
rect 258690 337958 258718 338028
rect 258678 337952 258730 337958
rect 258678 337894 258730 337900
rect 258782 337736 258810 338028
rect 258874 337958 258902 338028
rect 258966 337958 258994 338028
rect 258862 337952 258914 337958
rect 258862 337894 258914 337900
rect 258954 337952 259006 337958
rect 258954 337894 259006 337900
rect 259058 337770 259086 338028
rect 258598 337708 258672 337736
rect 258540 337544 258592 337550
rect 258540 337486 258592 337492
rect 258368 336382 258488 336410
rect 258262 336152 258318 336161
rect 258262 336087 258318 336096
rect 258078 336016 258134 336025
rect 258078 335951 258134 335960
rect 258170 335880 258226 335889
rect 258170 335815 258226 335824
rect 258184 335510 258212 335815
rect 258172 335504 258224 335510
rect 258172 335446 258224 335452
rect 258368 335442 258396 336382
rect 258448 336320 258500 336326
rect 258448 336262 258500 336268
rect 258356 335436 258408 335442
rect 258356 335378 258408 335384
rect 258460 332594 258488 336262
rect 258368 332566 258488 332594
rect 257988 326732 258040 326738
rect 257988 326674 258040 326680
rect 257988 326596 258040 326602
rect 257988 326538 258040 326544
rect 258000 97986 258028 326538
rect 258264 326392 258316 326398
rect 258264 326334 258316 326340
rect 257988 97980 258040 97986
rect 257988 97922 258040 97928
rect 257896 97776 257948 97782
rect 257896 97718 257948 97724
rect 257802 93936 257858 93945
rect 257802 93871 257858 93880
rect 257986 93800 258042 93809
rect 257986 93735 258042 93744
rect 258000 84289 258028 93735
rect 257986 84280 258042 84289
rect 257986 84215 258042 84224
rect 257986 84144 258042 84153
rect 257986 84079 258042 84088
rect 258000 74633 258028 84079
rect 257986 74624 258042 74633
rect 257986 74559 258042 74568
rect 257986 74488 258042 74497
rect 257986 74423 258042 74432
rect 258000 64977 258028 74423
rect 257986 64968 258042 64977
rect 257986 64903 258042 64912
rect 257986 64832 258042 64841
rect 257986 64767 258042 64776
rect 258000 55321 258028 64767
rect 257986 55312 258042 55321
rect 257986 55247 258042 55256
rect 257986 55176 258042 55185
rect 257986 55111 258042 55120
rect 258000 45665 258028 55111
rect 257986 45656 258042 45665
rect 257986 45591 258042 45600
rect 257986 45520 258042 45529
rect 257986 45455 258042 45464
rect 258000 36009 258028 45455
rect 257986 36000 258042 36009
rect 257986 35935 258042 35944
rect 257986 35864 258042 35873
rect 257986 35799 258042 35808
rect 258000 26353 258028 35799
rect 257986 26344 258042 26353
rect 257986 26279 258042 26288
rect 257986 26208 258042 26217
rect 257986 26143 258042 26152
rect 258000 16697 258028 26143
rect 257986 16688 258042 16697
rect 257986 16623 258042 16632
rect 257986 16552 258042 16561
rect 257986 16487 258042 16496
rect 258000 7041 258028 16487
rect 258276 7750 258304 326334
rect 258368 159390 258396 332566
rect 258552 332246 258580 337486
rect 258540 332240 258592 332246
rect 258540 332182 258592 332188
rect 258448 326188 258500 326194
rect 258448 326130 258500 326136
rect 258460 177886 258488 326130
rect 258540 323060 258592 323066
rect 258540 323002 258592 323008
rect 258448 177880 258500 177886
rect 258448 177822 258500 177828
rect 258356 159384 258408 159390
rect 258356 159326 258408 159332
rect 258446 158808 258502 158817
rect 258446 158743 258502 158752
rect 258264 7744 258316 7750
rect 258264 7686 258316 7692
rect 257986 7032 258042 7041
rect 257986 6967 258042 6976
rect 257712 3800 257764 3806
rect 257712 3742 257764 3748
rect 257528 3528 257580 3534
rect 257528 3470 257580 3476
rect 257436 3460 257488 3466
rect 257436 3402 257488 3408
rect 257038 354 257150 480
rect 256712 326 257150 354
rect 257038 -960 257150 326
rect 258234 354 258346 480
rect 258460 354 258488 158743
rect 258552 6390 258580 323002
rect 258644 321554 258672 337708
rect 258736 337708 258810 337736
rect 258920 337742 259086 337770
rect 258736 323066 258764 337708
rect 258816 337612 258868 337618
rect 258816 337554 258868 337560
rect 258828 334966 258856 337554
rect 258816 334960 258868 334966
rect 258816 334902 258868 334908
rect 258920 332594 258948 337742
rect 259150 337736 259178 338028
rect 259242 337958 259270 338028
rect 259334 337963 259362 338028
rect 259230 337952 259282 337958
rect 259230 337894 259282 337900
rect 259320 337954 259376 337963
rect 259426 337958 259454 338028
rect 259518 337958 259546 338028
rect 259610 337958 259638 338028
rect 259320 337889 259376 337898
rect 259414 337952 259466 337958
rect 259414 337894 259466 337900
rect 259506 337952 259558 337958
rect 259506 337894 259558 337900
rect 259598 337952 259650 337958
rect 259598 337894 259650 337900
rect 259702 337890 259730 338028
rect 259794 337963 259822 338028
rect 259780 337954 259836 337963
rect 259886 337958 259914 338028
rect 259978 337958 260006 338028
rect 259690 337884 259742 337890
rect 259780 337889 259836 337898
rect 259874 337952 259926 337958
rect 259874 337894 259926 337900
rect 259966 337952 260018 337958
rect 259966 337894 260018 337900
rect 259690 337826 259742 337832
rect 259460 337816 259512 337822
rect 259274 337784 259330 337793
rect 259150 337708 259224 337736
rect 259874 337816 259926 337822
rect 259460 337758 259512 337764
rect 259872 337784 259874 337793
rect 260070 337804 260098 338028
rect 260162 337929 260190 338028
rect 260254 337958 260282 338028
rect 260242 337952 260294 337958
rect 260148 337920 260204 337929
rect 260242 337894 260294 337900
rect 260148 337855 260204 337864
rect 259926 337784 259928 337793
rect 259274 337719 259330 337728
rect 259000 337612 259052 337618
rect 259000 337554 259052 337560
rect 259012 334422 259040 337554
rect 259196 336326 259224 337708
rect 259184 336320 259236 336326
rect 259184 336262 259236 336268
rect 259184 335980 259236 335986
rect 259184 335922 259236 335928
rect 259000 334416 259052 334422
rect 259000 334358 259052 334364
rect 258920 332566 259040 332594
rect 259012 326194 259040 332566
rect 259000 326188 259052 326194
rect 259000 326130 259052 326136
rect 258724 323060 258776 323066
rect 258724 323002 258776 323008
rect 259196 321554 259224 335922
rect 259288 326398 259316 337719
rect 259368 337680 259420 337686
rect 259368 337622 259420 337628
rect 259380 327894 259408 337622
rect 259472 335850 259500 337758
rect 259552 337748 259604 337754
rect 259872 337719 259928 337728
rect 259978 337776 260098 337804
rect 259978 337736 260006 337776
rect 260346 337736 260374 338028
rect 260438 337958 260466 338028
rect 260530 337958 260558 338028
rect 260426 337952 260478 337958
rect 260426 337894 260478 337900
rect 260518 337952 260570 337958
rect 260518 337894 260570 337900
rect 259978 337708 260052 337736
rect 259552 337690 259604 337696
rect 259460 335844 259512 335850
rect 259460 335786 259512 335792
rect 259564 335753 259592 337690
rect 259644 337544 259696 337550
rect 259644 337486 259696 337492
rect 259550 335744 259606 335753
rect 259550 335679 259606 335688
rect 259656 334529 259684 337486
rect 259828 337476 259880 337482
rect 259828 337418 259880 337424
rect 259736 336320 259788 336326
rect 259736 336262 259788 336268
rect 259642 334520 259698 334529
rect 259642 334455 259698 334464
rect 259748 332594 259776 336262
rect 259564 332566 259776 332594
rect 259564 330750 259592 332566
rect 259552 330744 259604 330750
rect 259552 330686 259604 330692
rect 259368 327888 259420 327894
rect 259368 327830 259420 327836
rect 259276 326392 259328 326398
rect 259276 326334 259328 326340
rect 259736 324216 259788 324222
rect 259736 324158 259788 324164
rect 258644 321526 258764 321554
rect 259196 321526 259408 321554
rect 258736 8090 258764 321526
rect 258998 158536 259054 158545
rect 258998 158471 259054 158480
rect 259012 97850 259040 158471
rect 259276 155916 259328 155922
rect 259276 155858 259328 155864
rect 259092 155848 259144 155854
rect 259092 155790 259144 155796
rect 259000 97844 259052 97850
rect 259000 97786 259052 97792
rect 258724 8084 258776 8090
rect 258724 8026 258776 8032
rect 258540 6384 258592 6390
rect 258540 6326 258592 6332
rect 259104 3398 259132 155790
rect 259184 155780 259236 155786
rect 259184 155722 259236 155728
rect 259196 4010 259224 155722
rect 259184 4004 259236 4010
rect 259184 3946 259236 3952
rect 259092 3392 259144 3398
rect 259092 3334 259144 3340
rect 259288 3262 259316 155858
rect 259380 3670 259408 321526
rect 259748 161474 259776 324158
rect 259472 161446 259776 161474
rect 259472 155378 259500 161446
rect 259552 161288 259604 161294
rect 259552 161230 259604 161236
rect 259460 155372 259512 155378
rect 259460 155314 259512 155320
rect 259564 97714 259592 161230
rect 259840 158030 259868 337418
rect 259920 337408 259972 337414
rect 259920 337350 259972 337356
rect 259932 335170 259960 337350
rect 260024 335918 260052 337708
rect 260300 337708 260374 337736
rect 260196 337680 260248 337686
rect 260102 337648 260158 337657
rect 260196 337622 260248 337628
rect 260102 337583 260158 337592
rect 260012 335912 260064 335918
rect 260012 335854 260064 335860
rect 259920 335164 259972 335170
rect 259920 335106 259972 335112
rect 259920 332240 259972 332246
rect 259920 332182 259972 332188
rect 259932 158030 259960 332182
rect 260012 326392 260064 326398
rect 260012 326334 260064 326340
rect 260116 326346 260144 337583
rect 260208 326482 260236 337622
rect 260300 336326 260328 337708
rect 260622 337668 260650 338028
rect 260714 337822 260742 338028
rect 260702 337816 260754 337822
rect 260702 337758 260754 337764
rect 260806 337736 260834 338028
rect 260898 337804 260926 338028
rect 260990 337929 261018 338028
rect 260976 337920 261032 337929
rect 260976 337855 261032 337864
rect 261082 337804 261110 338028
rect 261174 337890 261202 338028
rect 261266 337958 261294 338028
rect 261254 337952 261306 337958
rect 261254 337894 261306 337900
rect 261162 337884 261214 337890
rect 261162 337826 261214 337832
rect 260898 337776 260972 337804
rect 260806 337708 260880 337736
rect 260622 337640 260788 337668
rect 260564 337544 260616 337550
rect 260564 337486 260616 337492
rect 260472 337476 260524 337482
rect 260472 337418 260524 337424
rect 260288 336320 260340 336326
rect 260288 336262 260340 336268
rect 260288 335912 260340 335918
rect 260288 335854 260340 335860
rect 260300 330614 260328 335854
rect 260288 330608 260340 330614
rect 260288 330550 260340 330556
rect 260208 326454 260420 326482
rect 259828 158024 259880 158030
rect 259828 157966 259880 157972
rect 259920 158024 259972 158030
rect 259920 157966 259972 157972
rect 259828 157480 259880 157486
rect 259828 157422 259880 157428
rect 259644 156732 259696 156738
rect 259644 156674 259696 156680
rect 259552 97708 259604 97714
rect 259552 97650 259604 97656
rect 259656 6914 259684 156674
rect 259736 156664 259788 156670
rect 259736 156606 259788 156612
rect 259748 100502 259776 156606
rect 259736 100496 259788 100502
rect 259736 100438 259788 100444
rect 259840 16574 259868 157422
rect 259920 156052 259972 156058
rect 259920 155994 259972 156000
rect 259932 155242 259960 155994
rect 260024 155446 260052 326334
rect 260116 326318 260328 326346
rect 260196 326256 260248 326262
rect 260196 326198 260248 326204
rect 260208 320890 260236 326198
rect 260196 320884 260248 320890
rect 260196 320826 260248 320832
rect 260300 171134 260328 326318
rect 260392 326262 260420 326454
rect 260380 326256 260432 326262
rect 260380 326198 260432 326204
rect 260300 171106 260420 171134
rect 260392 156058 260420 171106
rect 260380 156052 260432 156058
rect 260380 155994 260432 156000
rect 260288 155712 260340 155718
rect 260286 155680 260288 155689
rect 260340 155680 260342 155689
rect 260286 155615 260342 155624
rect 260484 155446 260512 337418
rect 260576 324222 260604 337486
rect 260656 337476 260708 337482
rect 260656 337418 260708 337424
rect 260668 326398 260696 337418
rect 260760 332382 260788 337640
rect 260852 335374 260880 337708
rect 260944 336666 260972 337776
rect 261036 337776 261110 337804
rect 260932 336660 260984 336666
rect 260932 336602 260984 336608
rect 260840 335368 260892 335374
rect 261036 335345 261064 337776
rect 261208 337748 261260 337754
rect 261208 337690 261260 337696
rect 261220 337657 261248 337690
rect 261358 337668 261386 338028
rect 261450 337770 261478 338028
rect 261542 337963 261570 338028
rect 261528 337954 261584 337963
rect 261634 337958 261662 338028
rect 261726 337958 261754 338028
rect 261528 337889 261584 337898
rect 261622 337952 261674 337958
rect 261622 337894 261674 337900
rect 261714 337952 261766 337958
rect 261714 337894 261766 337900
rect 261818 337804 261846 338028
rect 261772 337776 261846 337804
rect 261450 337742 261616 337770
rect 261206 337648 261262 337657
rect 261116 337612 261168 337618
rect 261358 337640 261432 337668
rect 261206 337583 261262 337592
rect 261116 337554 261168 337560
rect 260840 335310 260892 335316
rect 261022 335336 261078 335345
rect 261022 335271 261078 335280
rect 260748 332376 260800 332382
rect 260748 332318 260800 332324
rect 260748 331288 260800 331294
rect 260748 331230 260800 331236
rect 260656 326392 260708 326398
rect 260656 326334 260708 326340
rect 260564 324216 260616 324222
rect 260564 324158 260616 324164
rect 260564 158024 260616 158030
rect 260564 157966 260616 157972
rect 260576 155938 260604 157966
rect 260760 156670 260788 331230
rect 261024 323060 261076 323066
rect 261024 323002 261076 323008
rect 261036 156806 261064 323002
rect 261128 158098 261156 337554
rect 261208 337544 261260 337550
rect 261208 337486 261260 337492
rect 261220 333810 261248 337486
rect 261300 335776 261352 335782
rect 261300 335718 261352 335724
rect 261208 333804 261260 333810
rect 261208 333746 261260 333752
rect 261312 332594 261340 335718
rect 261220 332566 261340 332594
rect 261220 331214 261248 332566
rect 261220 331186 261340 331214
rect 261312 330818 261340 331186
rect 261300 330812 261352 330818
rect 261300 330754 261352 330760
rect 261404 326602 261432 337640
rect 261482 337512 261538 337521
rect 261482 337447 261538 337456
rect 261392 326596 261444 326602
rect 261392 326538 261444 326544
rect 261496 326482 261524 337447
rect 261588 335782 261616 337742
rect 261668 337680 261720 337686
rect 261668 337622 261720 337628
rect 261576 335776 261628 335782
rect 261576 335718 261628 335724
rect 261576 335572 261628 335578
rect 261576 335514 261628 335520
rect 261220 326454 261524 326482
rect 261220 158166 261248 326454
rect 261300 326392 261352 326398
rect 261588 326346 261616 335514
rect 261300 326334 261352 326340
rect 261312 159458 261340 326334
rect 261392 326324 261444 326330
rect 261392 326266 261444 326272
rect 261496 326318 261616 326346
rect 261404 160721 261432 326266
rect 261390 160712 261446 160721
rect 261390 160647 261446 160656
rect 261300 159452 261352 159458
rect 261300 159394 261352 159400
rect 261208 158160 261260 158166
rect 261208 158102 261260 158108
rect 261116 158092 261168 158098
rect 261116 158034 261168 158040
rect 261496 157826 261524 326318
rect 261680 321554 261708 337622
rect 261772 335714 261800 337776
rect 261910 337736 261938 338028
rect 262002 337963 262030 338028
rect 261988 337954 262044 337963
rect 262094 337958 262122 338028
rect 261988 337889 262044 337898
rect 262082 337952 262134 337958
rect 262082 337894 262134 337900
rect 262186 337890 262214 338028
rect 262278 337958 262306 338028
rect 262266 337952 262318 337958
rect 262266 337894 262318 337900
rect 262174 337884 262226 337890
rect 262174 337826 262226 337832
rect 262036 337816 262088 337822
rect 262370 337793 262398 338028
rect 262462 337822 262490 338028
rect 262450 337816 262502 337822
rect 262036 337758 262088 337764
rect 262356 337784 262412 337793
rect 261864 337708 261938 337736
rect 261760 335708 261812 335714
rect 261760 335650 261812 335656
rect 261760 326596 261812 326602
rect 261760 326538 261812 326544
rect 261588 321526 261708 321554
rect 261484 157820 261536 157826
rect 261484 157762 261536 157768
rect 261024 156800 261076 156806
rect 261024 156742 261076 156748
rect 260748 156664 260800 156670
rect 260748 156606 260800 156612
rect 260576 155910 260682 155938
rect 261588 155718 261616 321526
rect 261772 316034 261800 326538
rect 261864 326398 261892 337708
rect 261944 337612 261996 337618
rect 261944 337554 261996 337560
rect 261956 326534 261984 337554
rect 261944 326528 261996 326534
rect 261944 326470 261996 326476
rect 261852 326392 261904 326398
rect 261852 326334 261904 326340
rect 262048 326330 262076 337758
rect 262220 337748 262272 337754
rect 262450 337758 262502 337764
rect 262554 337770 262582 338028
rect 262646 337963 262674 338028
rect 262632 337954 262688 337963
rect 262738 337958 262766 338028
rect 262632 337889 262688 337898
rect 262726 337952 262778 337958
rect 262830 337929 262858 338028
rect 262922 337958 262950 338028
rect 263014 337958 263042 338028
rect 263106 337958 263134 338028
rect 263198 337963 263226 338028
rect 262910 337952 262962 337958
rect 262726 337894 262778 337900
rect 262816 337920 262872 337929
rect 262910 337894 262962 337900
rect 263002 337952 263054 337958
rect 263002 337894 263054 337900
rect 263094 337952 263146 337958
rect 263094 337894 263146 337900
rect 263184 337954 263240 337963
rect 263184 337889 263240 337898
rect 262816 337855 262872 337864
rect 263290 337822 263318 338028
rect 262956 337816 263008 337822
rect 262554 337742 262674 337770
rect 263278 337816 263330 337822
rect 262956 337758 263008 337764
rect 263046 337784 263102 337793
rect 262356 337719 262412 337728
rect 262646 337736 262674 337742
rect 262646 337708 262720 337736
rect 262220 337690 262272 337696
rect 262126 337648 262182 337657
rect 262126 337583 262182 337592
rect 262036 326324 262088 326330
rect 262036 326266 262088 326272
rect 262140 323066 262168 337583
rect 262232 337142 262260 337690
rect 262310 337648 262366 337657
rect 262310 337583 262366 337592
rect 262588 337612 262640 337618
rect 262220 337136 262272 337142
rect 262220 337078 262272 337084
rect 262324 336530 262352 337583
rect 262588 337554 262640 337560
rect 262496 337544 262548 337550
rect 262496 337486 262548 337492
rect 262312 336524 262364 336530
rect 262312 336466 262364 336472
rect 262508 331214 262536 337486
rect 262600 336002 262628 337554
rect 262692 336258 262720 337708
rect 262680 336252 262732 336258
rect 262680 336194 262732 336200
rect 262600 335974 262904 336002
rect 262680 335912 262732 335918
rect 262586 335880 262642 335889
rect 262680 335854 262732 335860
rect 262586 335815 262642 335824
rect 262416 331186 262536 331214
rect 262128 323060 262180 323066
rect 262128 323002 262180 323008
rect 261680 316006 261800 316034
rect 261680 156602 261708 316006
rect 262416 159594 262444 331186
rect 262496 326460 262548 326466
rect 262496 326402 262548 326408
rect 262508 159662 262536 326402
rect 262496 159656 262548 159662
rect 262496 159598 262548 159604
rect 262404 159588 262456 159594
rect 262404 159530 262456 159536
rect 262600 159526 262628 335815
rect 262692 332314 262720 335854
rect 262680 332308 262732 332314
rect 262680 332250 262732 332256
rect 262680 326392 262732 326398
rect 262680 326334 262732 326340
rect 262588 159520 262640 159526
rect 262588 159462 262640 159468
rect 262692 156874 262720 326334
rect 262876 158234 262904 335974
rect 262968 335918 262996 337758
rect 263278 337758 263330 337764
rect 263046 337719 263102 337728
rect 262956 335912 263008 335918
rect 262956 335854 263008 335860
rect 263060 335034 263088 337719
rect 263140 337680 263192 337686
rect 263382 337668 263410 338028
rect 263140 337622 263192 337628
rect 263336 337640 263410 337668
rect 263152 337210 263180 337622
rect 263232 337476 263284 337482
rect 263232 337418 263284 337424
rect 263140 337204 263192 337210
rect 263140 337146 263192 337152
rect 263048 335028 263100 335034
rect 263048 334970 263100 334976
rect 263244 326466 263272 337418
rect 263232 326460 263284 326466
rect 263232 326402 263284 326408
rect 263336 326398 263364 337640
rect 263474 337600 263502 338028
rect 263566 337958 263594 338028
rect 263658 337958 263686 338028
rect 263554 337952 263606 337958
rect 263554 337894 263606 337900
rect 263646 337952 263698 337958
rect 263646 337894 263698 337900
rect 263750 337793 263778 338028
rect 263842 337890 263870 338028
rect 263934 337929 263962 338028
rect 264026 337958 264054 338028
rect 264014 337952 264066 337958
rect 263920 337920 263976 337929
rect 263830 337884 263882 337890
rect 264014 337894 264066 337900
rect 263920 337855 263976 337864
rect 263830 337826 263882 337832
rect 263736 337784 263792 337793
rect 264118 337770 264146 338028
rect 264210 337822 264238 338028
rect 263736 337719 263792 337728
rect 263876 337748 263928 337754
rect 263876 337690 263928 337696
rect 263980 337742 264146 337770
rect 264198 337816 264250 337822
rect 264198 337758 264250 337764
rect 263428 337572 263502 337600
rect 263428 335102 263456 337572
rect 263508 337476 263560 337482
rect 263508 337418 263560 337424
rect 263692 337476 263744 337482
rect 263692 337418 263744 337424
rect 263416 335096 263468 335102
rect 263416 335038 263468 335044
rect 263520 331214 263548 337418
rect 263704 336802 263732 337418
rect 263692 336796 263744 336802
rect 263692 336738 263744 336744
rect 263888 336705 263916 337690
rect 263874 336696 263930 336705
rect 263874 336631 263930 336640
rect 263980 333810 264008 337742
rect 264060 337680 264112 337686
rect 264302 337668 264330 338028
rect 264394 337822 264422 338028
rect 264486 337929 264514 338028
rect 264472 337920 264528 337929
rect 264472 337855 264528 337864
rect 264382 337816 264434 337822
rect 264382 337758 264434 337764
rect 264060 337622 264112 337628
rect 264256 337640 264330 337668
rect 264428 337680 264480 337686
rect 263968 333804 264020 333810
rect 263968 333746 264020 333752
rect 263428 331186 263548 331214
rect 263428 330886 263456 331186
rect 263506 331120 263562 331129
rect 263506 331055 263562 331064
rect 263416 330880 263468 330886
rect 263416 330822 263468 330828
rect 263324 326392 263376 326398
rect 263324 326334 263376 326340
rect 263520 321609 263548 331055
rect 263784 330676 263836 330682
rect 263784 330618 263836 330624
rect 263506 321600 263562 321609
rect 263506 321535 263562 321544
rect 263796 158302 263824 330618
rect 263968 330608 264020 330614
rect 263968 330550 264020 330556
rect 263876 330472 263928 330478
rect 263876 330414 263928 330420
rect 263888 159730 263916 330414
rect 263980 159866 264008 330550
rect 264072 330546 264100 337622
rect 264256 337600 264284 337640
rect 264578 337668 264606 338028
rect 264670 337890 264698 338028
rect 264762 337890 264790 338028
rect 264658 337884 264710 337890
rect 264658 337826 264710 337832
rect 264750 337884 264802 337890
rect 264750 337826 264802 337832
rect 264702 337784 264758 337793
rect 264854 337770 264882 338028
rect 264702 337719 264758 337728
rect 264808 337742 264882 337770
rect 264428 337622 264480 337628
rect 264532 337640 264606 337668
rect 264256 337572 264330 337600
rect 264302 337532 264330 337572
rect 264302 337504 264376 337532
rect 264244 337408 264296 337414
rect 264244 337350 264296 337356
rect 264152 337340 264204 337346
rect 264152 337282 264204 337288
rect 264060 330540 264112 330546
rect 264060 330482 264112 330488
rect 264060 330404 264112 330410
rect 264060 330346 264112 330352
rect 263968 159860 264020 159866
rect 263968 159802 264020 159808
rect 264072 159798 264100 330346
rect 264164 160546 264192 337282
rect 264256 336190 264284 337350
rect 264244 336184 264296 336190
rect 264244 336126 264296 336132
rect 264244 334620 264296 334626
rect 264244 334562 264296 334568
rect 264152 160540 264204 160546
rect 264152 160482 264204 160488
rect 264060 159792 264112 159798
rect 264060 159734 264112 159740
rect 263876 159724 263928 159730
rect 263876 159666 263928 159672
rect 263784 158296 263836 158302
rect 263784 158238 263836 158244
rect 262864 158228 262916 158234
rect 262864 158170 262916 158176
rect 264256 157078 264284 334562
rect 264348 330682 264376 337504
rect 264336 330676 264388 330682
rect 264336 330618 264388 330624
rect 264336 330540 264388 330546
rect 264336 330482 264388 330488
rect 264244 157072 264296 157078
rect 264244 157014 264296 157020
rect 264348 157010 264376 330482
rect 264440 330478 264468 337622
rect 264428 330472 264480 330478
rect 264428 330414 264480 330420
rect 264532 330410 264560 337640
rect 264612 337544 264664 337550
rect 264612 337486 264664 337492
rect 264624 334626 264652 337486
rect 264612 334620 264664 334626
rect 264612 334562 264664 334568
rect 264716 331214 264744 337719
rect 264624 331186 264744 331214
rect 264520 330404 264572 330410
rect 264520 330346 264572 330352
rect 264624 330342 264652 331186
rect 264808 330614 264836 337742
rect 264946 337668 264974 338028
rect 265038 337890 265066 338028
rect 265130 337963 265158 338028
rect 265116 337954 265172 337963
rect 265026 337884 265078 337890
rect 265116 337889 265172 337898
rect 265026 337826 265078 337832
rect 265072 337748 265124 337754
rect 265072 337690 265124 337696
rect 264900 337640 264974 337668
rect 264900 330750 264928 337640
rect 264980 337476 265032 337482
rect 264980 337418 265032 337424
rect 264992 336598 265020 337418
rect 264980 336592 265032 336598
rect 264980 336534 265032 336540
rect 265084 335481 265112 337690
rect 265222 337668 265250 338028
rect 265314 337890 265342 338028
rect 265406 337929 265434 338028
rect 265498 337958 265526 338028
rect 265590 337963 265618 338028
rect 265486 337952 265538 337958
rect 265392 337920 265448 337929
rect 265302 337884 265354 337890
rect 265486 337894 265538 337900
rect 265576 337954 265632 337963
rect 265576 337889 265632 337898
rect 265682 337890 265710 338028
rect 265392 337855 265448 337864
rect 265670 337884 265722 337890
rect 265302 337826 265354 337832
rect 265670 337826 265722 337832
rect 265438 337784 265494 337793
rect 265348 337748 265400 337754
rect 265774 337770 265802 338028
rect 265728 337754 265802 337770
rect 265438 337719 265494 337728
rect 265716 337748 265802 337754
rect 265348 337690 265400 337696
rect 265222 337640 265296 337668
rect 265164 337544 265216 337550
rect 265164 337486 265216 337492
rect 265070 335472 265126 335481
rect 265070 335407 265126 335416
rect 264888 330744 264940 330750
rect 264888 330686 264940 330692
rect 264796 330608 264848 330614
rect 264796 330550 264848 330556
rect 264612 330336 264664 330342
rect 264612 330278 264664 330284
rect 264520 158364 264572 158370
rect 264520 158306 264572 158312
rect 264336 157004 264388 157010
rect 264336 156946 264388 156952
rect 262680 156868 262732 156874
rect 262680 156810 262732 156816
rect 261668 156596 261720 156602
rect 261668 156538 261720 156544
rect 264532 155924 264560 158306
rect 265176 156738 265204 337486
rect 265268 335617 265296 337640
rect 265254 335608 265310 335617
rect 265360 335578 265388 337690
rect 265254 335543 265310 335552
rect 265348 335572 265400 335578
rect 265348 335514 265400 335520
rect 265452 335481 265480 337719
rect 265768 337742 265802 337748
rect 265866 337770 265894 338028
rect 265958 337890 265986 338028
rect 265946 337884 265998 337890
rect 265946 337826 265998 337832
rect 266050 337770 266078 338028
rect 266142 337895 266170 338028
rect 266128 337886 266184 337895
rect 266128 337821 266184 337830
rect 265866 337742 265940 337770
rect 266050 337742 266124 337770
rect 265716 337690 265768 337696
rect 265624 337680 265676 337686
rect 265530 337648 265586 337657
rect 265624 337622 265676 337628
rect 265530 337583 265586 337592
rect 265438 335472 265494 335481
rect 265438 335407 265494 335416
rect 265440 334620 265492 334626
rect 265440 334562 265492 334568
rect 265256 330540 265308 330546
rect 265256 330482 265308 330488
rect 265268 157486 265296 330482
rect 265348 329724 265400 329730
rect 265348 329666 265400 329672
rect 265360 158642 265388 329666
rect 265452 160682 265480 334562
rect 265544 330546 265572 337583
rect 265636 333470 265664 337622
rect 265716 337612 265768 337618
rect 265912 337600 265940 337742
rect 266096 337618 266124 337742
rect 266234 337668 266262 338028
rect 266188 337640 266262 337668
rect 266084 337612 266136 337618
rect 265912 337572 266032 337600
rect 265716 337554 265768 337560
rect 265728 334370 265756 337554
rect 265900 337476 265952 337482
rect 265900 337418 265952 337424
rect 265808 337408 265860 337414
rect 265808 337350 265860 337356
rect 265820 334626 265848 337350
rect 265808 334620 265860 334626
rect 265808 334562 265860 334568
rect 265728 334342 265848 334370
rect 265716 334280 265768 334286
rect 265716 334222 265768 334228
rect 265624 333464 265676 333470
rect 265624 333406 265676 333412
rect 265532 330540 265584 330546
rect 265532 330482 265584 330488
rect 265532 330404 265584 330410
rect 265532 330346 265584 330352
rect 265440 160676 265492 160682
rect 265440 160618 265492 160624
rect 265348 158636 265400 158642
rect 265348 158578 265400 158584
rect 265256 157480 265308 157486
rect 265256 157422 265308 157428
rect 265164 156732 265216 156738
rect 265164 156674 265216 156680
rect 265544 155922 265572 330346
rect 265728 316034 265756 334222
rect 265820 332994 265848 334342
rect 265808 332988 265860 332994
rect 265808 332930 265860 332936
rect 265912 316034 265940 337418
rect 266004 331294 266032 337572
rect 266084 337554 266136 337560
rect 266082 337512 266138 337521
rect 266082 337447 266138 337456
rect 265992 331288 266044 331294
rect 265992 331230 266044 331236
rect 266096 330410 266124 337447
rect 266084 330404 266136 330410
rect 266084 330346 266136 330352
rect 266188 329730 266216 337640
rect 266326 337532 266354 338028
rect 266418 337770 266446 338028
rect 266510 337890 266538 338028
rect 266602 337890 266630 338028
rect 266694 337929 266722 338028
rect 266680 337920 266736 337929
rect 266498 337884 266550 337890
rect 266498 337826 266550 337832
rect 266590 337884 266642 337890
rect 266680 337855 266736 337864
rect 266590 337826 266642 337832
rect 266418 337742 266492 337770
rect 266280 337504 266354 337532
rect 266280 336258 266308 337504
rect 266358 336832 266414 336841
rect 266358 336767 266414 336776
rect 266268 336252 266320 336258
rect 266268 336194 266320 336200
rect 266372 336138 266400 336767
rect 266280 336110 266400 336138
rect 266280 334286 266308 336110
rect 266268 334280 266320 334286
rect 266268 334222 266320 334228
rect 266464 330818 266492 337742
rect 266636 337748 266688 337754
rect 266786 337736 266814 338028
rect 266878 337804 266906 338028
rect 266970 337958 266998 338028
rect 267062 337958 267090 338028
rect 267154 337958 267182 338028
rect 266958 337952 267010 337958
rect 266958 337894 267010 337900
rect 267050 337952 267102 337958
rect 267050 337894 267102 337900
rect 267142 337952 267194 337958
rect 267142 337894 267194 337900
rect 267246 337890 267274 338028
rect 267338 337890 267366 338028
rect 267234 337884 267286 337890
rect 267234 337826 267286 337832
rect 267326 337884 267378 337890
rect 267326 337826 267378 337832
rect 267004 337816 267056 337822
rect 266878 337776 266952 337804
rect 266786 337708 266860 337736
rect 266636 337690 266688 337696
rect 266542 337648 266598 337657
rect 266648 337634 266676 337690
rect 266648 337606 266768 337634
rect 266542 337583 266598 337592
rect 266452 330812 266504 330818
rect 266452 330754 266504 330760
rect 266556 330698 266584 337583
rect 266636 337544 266688 337550
rect 266636 337486 266688 337492
rect 266464 330670 266584 330698
rect 266176 329724 266228 329730
rect 266176 329666 266228 329672
rect 265636 316006 265756 316034
rect 265820 316006 265940 316034
rect 265636 158370 265664 316006
rect 265624 158364 265676 158370
rect 265624 158306 265676 158312
rect 265532 155916 265584 155922
rect 265532 155858 265584 155864
rect 261576 155712 261628 155718
rect 261576 155654 261628 155660
rect 265820 155514 265848 316006
rect 266464 155689 266492 330670
rect 266544 330608 266596 330614
rect 266544 330550 266596 330556
rect 266556 155854 266584 330550
rect 266648 157962 266676 337486
rect 266740 334626 266768 337606
rect 266728 334620 266780 334626
rect 266728 334562 266780 334568
rect 266728 330404 266780 330410
rect 266728 330346 266780 330352
rect 266740 158438 266768 330346
rect 266832 158574 266860 337708
rect 266924 330682 266952 337776
rect 267430 337770 267458 338028
rect 267522 337958 267550 338028
rect 267510 337952 267562 337958
rect 267614 337929 267642 338028
rect 267510 337894 267562 337900
rect 267600 337920 267656 337929
rect 267600 337855 267656 337864
rect 267004 337758 267056 337764
rect 266912 330676 266964 330682
rect 266912 330618 266964 330624
rect 267016 330562 267044 337758
rect 267096 337748 267148 337754
rect 267096 337690 267148 337696
rect 267292 337742 267458 337770
rect 266924 330534 267044 330562
rect 266820 158568 266872 158574
rect 266820 158510 266872 158516
rect 266728 158432 266780 158438
rect 266728 158374 266780 158380
rect 266924 158302 266952 330534
rect 267004 330472 267056 330478
rect 267004 330414 267056 330420
rect 267016 161430 267044 330414
rect 267004 161424 267056 161430
rect 267004 161366 267056 161372
rect 267108 161090 267136 337690
rect 267188 337680 267240 337686
rect 267188 337622 267240 337628
rect 267200 335354 267228 337622
rect 267292 336938 267320 337742
rect 267464 337680 267516 337686
rect 267706 337668 267734 338028
rect 267464 337622 267516 337628
rect 267660 337640 267734 337668
rect 267372 337612 267424 337618
rect 267372 337554 267424 337560
rect 267280 336932 267332 336938
rect 267280 336874 267332 336880
rect 267200 335326 267320 335354
rect 267188 334620 267240 334626
rect 267188 334562 267240 334568
rect 267200 161226 267228 334562
rect 267292 325694 267320 335326
rect 267384 330410 267412 337554
rect 267476 336705 267504 337622
rect 267462 336696 267518 336705
rect 267462 336631 267518 336640
rect 267660 335354 267688 337640
rect 267798 337634 267826 338028
rect 267890 337770 267918 338028
rect 267982 337929 268010 338028
rect 268074 337958 268102 338028
rect 268062 337952 268114 337958
rect 267968 337920 268024 337929
rect 268062 337894 268114 337900
rect 267968 337855 268024 337864
rect 268014 337784 268070 337793
rect 267890 337742 267964 337770
rect 267798 337606 267872 337634
rect 267740 337544 267792 337550
rect 267740 337486 267792 337492
rect 267752 336122 267780 337486
rect 267740 336116 267792 336122
rect 267740 336058 267792 336064
rect 267660 335326 267780 335354
rect 267372 330404 267424 330410
rect 267372 330346 267424 330352
rect 267752 330274 267780 335326
rect 267740 330268 267792 330274
rect 267740 330210 267792 330216
rect 267292 325666 267596 325694
rect 267188 161220 267240 161226
rect 267188 161162 267240 161168
rect 267096 161084 267148 161090
rect 267096 161026 267148 161032
rect 266912 158296 266964 158302
rect 266912 158238 266964 158244
rect 266636 157956 266688 157962
rect 266636 157898 266688 157904
rect 266544 155848 266596 155854
rect 266544 155790 266596 155796
rect 267568 155786 267596 325666
rect 267556 155780 267608 155786
rect 267556 155722 267608 155728
rect 266450 155680 266506 155689
rect 267844 155650 267872 337606
rect 267936 158506 267964 337742
rect 268014 337719 268070 337728
rect 268028 330562 268056 337719
rect 268166 337634 268194 338028
rect 268258 337770 268286 338028
rect 268350 337890 268378 338028
rect 268338 337884 268390 337890
rect 268338 337826 268390 337832
rect 268442 337770 268470 338028
rect 268258 337742 268332 337770
rect 268166 337606 268240 337634
rect 268108 337476 268160 337482
rect 268108 337418 268160 337424
rect 268120 331214 268148 337418
rect 268212 336734 268240 337606
rect 268200 336728 268252 336734
rect 268200 336670 268252 336676
rect 268120 331186 268240 331214
rect 268028 330534 268148 330562
rect 268016 330472 268068 330478
rect 268016 330414 268068 330420
rect 268028 161022 268056 330414
rect 268016 161016 268068 161022
rect 268016 160958 268068 160964
rect 268120 160886 268148 330534
rect 268212 330478 268240 331186
rect 268304 330546 268332 337742
rect 268396 337742 268470 337770
rect 268292 330540 268344 330546
rect 268292 330482 268344 330488
rect 268200 330472 268252 330478
rect 268200 330414 268252 330420
rect 268292 330404 268344 330410
rect 268292 330346 268344 330352
rect 268200 330336 268252 330342
rect 268200 330278 268252 330284
rect 268108 160880 268160 160886
rect 268108 160822 268160 160828
rect 268212 160614 268240 330278
rect 268304 160954 268332 330346
rect 268292 160948 268344 160954
rect 268292 160890 268344 160896
rect 268396 160750 268424 337742
rect 268534 337668 268562 338028
rect 268626 337770 268654 338028
rect 268718 337929 268746 338028
rect 268704 337920 268760 337929
rect 268810 337890 268838 338028
rect 268704 337855 268760 337864
rect 268798 337884 268850 337890
rect 268798 337826 268850 337832
rect 268750 337784 268806 337793
rect 268626 337742 268700 337770
rect 268534 337640 268608 337668
rect 268476 337544 268528 337550
rect 268476 337486 268528 337492
rect 268488 335986 268516 337486
rect 268476 335980 268528 335986
rect 268476 335922 268528 335928
rect 268476 330540 268528 330546
rect 268476 330482 268528 330488
rect 268488 160818 268516 330482
rect 268580 330410 268608 337640
rect 268568 330404 268620 330410
rect 268568 330346 268620 330352
rect 268568 330268 268620 330274
rect 268568 330210 268620 330216
rect 268580 161158 268608 330210
rect 268568 161152 268620 161158
rect 268568 161094 268620 161100
rect 268476 160812 268528 160818
rect 268476 160754 268528 160760
rect 268384 160744 268436 160750
rect 268384 160686 268436 160692
rect 268200 160608 268252 160614
rect 268200 160550 268252 160556
rect 267924 158500 267976 158506
rect 267924 158442 267976 158448
rect 266450 155615 266506 155624
rect 267832 155644 267884 155650
rect 267832 155586 267884 155592
rect 268672 155582 268700 337742
rect 268902 337770 268930 338028
rect 268750 337719 268806 337728
rect 268856 337742 268930 337770
rect 268994 337770 269022 338028
rect 269086 337958 269114 338028
rect 269074 337952 269126 337958
rect 269074 337894 269126 337900
rect 269178 337890 269206 338028
rect 269166 337884 269218 337890
rect 269166 337826 269218 337832
rect 269270 337770 269298 338028
rect 269362 337958 269390 338028
rect 269350 337952 269402 337958
rect 269350 337894 269402 337900
rect 269454 337770 269482 338028
rect 269546 337822 269574 338028
rect 268994 337742 269068 337770
rect 268764 330342 268792 337719
rect 268856 335617 268884 337742
rect 268936 337680 268988 337686
rect 268936 337622 268988 337628
rect 268842 335608 268898 335617
rect 268842 335543 268898 335552
rect 268948 335481 268976 337622
rect 269040 335753 269068 337742
rect 269132 337742 269298 337770
rect 269408 337742 269482 337770
rect 269534 337816 269586 337822
rect 269534 337758 269586 337764
rect 269638 337770 269666 338028
rect 269730 337958 269758 338028
rect 269822 337958 269850 338028
rect 269718 337952 269770 337958
rect 269718 337894 269770 337900
rect 269810 337952 269862 337958
rect 269810 337894 269862 337900
rect 269764 337816 269816 337822
rect 269638 337742 269712 337770
rect 269914 337770 269942 338028
rect 269764 337758 269816 337764
rect 269026 335744 269082 335753
rect 269026 335679 269082 335688
rect 268934 335472 268990 335481
rect 268934 335407 268990 335416
rect 269132 330818 269160 337742
rect 269304 337680 269356 337686
rect 269304 337622 269356 337628
rect 269212 337544 269264 337550
rect 269212 337486 269264 337492
rect 269120 330812 269172 330818
rect 269120 330754 269172 330760
rect 269120 330676 269172 330682
rect 269120 330618 269172 330624
rect 268752 330336 268804 330342
rect 268752 330278 268804 330284
rect 269026 158672 269082 158681
rect 269026 158607 269082 158616
rect 269040 155924 269068 158607
rect 269132 155650 269160 330618
rect 269224 330562 269252 337486
rect 269316 330750 269344 337622
rect 269304 330744 269356 330750
rect 269304 330686 269356 330692
rect 269224 330534 269344 330562
rect 269212 330472 269264 330478
rect 269212 330414 269264 330420
rect 269224 155802 269252 330414
rect 269316 155938 269344 330534
rect 269408 330478 269436 337742
rect 269488 337680 269540 337686
rect 269488 337622 269540 337628
rect 269580 337680 269632 337686
rect 269580 337622 269632 337628
rect 269500 335481 269528 337622
rect 269486 335472 269542 335481
rect 269486 335407 269542 335416
rect 269592 330682 269620 337622
rect 269580 330676 269632 330682
rect 269580 330618 269632 330624
rect 269580 330540 269632 330546
rect 269580 330482 269632 330488
rect 269396 330472 269448 330478
rect 269396 330414 269448 330420
rect 269488 330472 269540 330478
rect 269488 330414 269540 330420
rect 269396 330336 269448 330342
rect 269396 330278 269448 330284
rect 269408 158710 269436 330278
rect 269396 158704 269448 158710
rect 269396 158646 269448 158652
rect 269500 158302 269528 330414
rect 269592 161401 269620 330482
rect 269578 161392 269634 161401
rect 269578 161327 269634 161336
rect 269684 160857 269712 337742
rect 269670 160848 269726 160857
rect 269670 160783 269726 160792
rect 269776 160585 269804 337758
rect 269868 337742 269942 337770
rect 269868 330546 269896 337742
rect 270006 337736 270034 338028
rect 270098 337890 270126 338028
rect 270086 337884 270138 337890
rect 270086 337826 270138 337832
rect 270190 337804 270218 338028
rect 270282 337958 270310 338028
rect 270374 337958 270402 338028
rect 270270 337952 270322 337958
rect 270270 337894 270322 337900
rect 270362 337952 270414 337958
rect 270466 337929 270494 338028
rect 270362 337894 270414 337900
rect 270452 337920 270508 337929
rect 270452 337855 270508 337864
rect 270408 337816 270460 337822
rect 270190 337776 270264 337804
rect 270006 337708 270172 337736
rect 270040 337612 270092 337618
rect 270040 337554 270092 337560
rect 270052 337006 270080 337554
rect 270040 337000 270092 337006
rect 270040 336942 270092 336948
rect 269948 335980 270000 335986
rect 269948 335922 270000 335928
rect 269856 330540 269908 330546
rect 269856 330482 269908 330488
rect 269960 330478 269988 335922
rect 270040 330744 270092 330750
rect 270040 330686 270092 330692
rect 269948 330472 270000 330478
rect 269948 330414 270000 330420
rect 270052 330290 270080 330686
rect 270144 330342 270172 337708
rect 270236 335986 270264 337776
rect 270406 337784 270408 337793
rect 270460 337784 270462 337793
rect 270558 337736 270586 338028
rect 270406 337719 270462 337728
rect 270512 337708 270586 337736
rect 270512 337634 270540 337708
rect 270650 337668 270678 338028
rect 270742 337958 270770 338028
rect 270834 337963 270862 338028
rect 270730 337952 270782 337958
rect 270730 337894 270782 337900
rect 270820 337954 270876 337963
rect 270820 337889 270876 337898
rect 270926 337890 270954 338028
rect 270914 337884 270966 337890
rect 270914 337826 270966 337832
rect 271018 337804 271046 338028
rect 271110 337958 271138 338028
rect 271202 337958 271230 338028
rect 271098 337952 271150 337958
rect 271098 337894 271150 337900
rect 271190 337952 271242 337958
rect 271190 337894 271242 337900
rect 271018 337776 271092 337804
rect 271294 337793 271322 338028
rect 271064 337770 271092 337776
rect 271280 337784 271336 337793
rect 271064 337742 271138 337770
rect 271110 337668 271138 337742
rect 271280 337719 271336 337728
rect 270650 337640 270724 337668
rect 270420 337606 270540 337634
rect 270420 336258 270448 337606
rect 270592 337544 270644 337550
rect 270592 337486 270644 337492
rect 270408 336252 270460 336258
rect 270408 336194 270460 336200
rect 270224 335980 270276 335986
rect 270224 335922 270276 335928
rect 270224 330812 270276 330818
rect 270224 330754 270276 330760
rect 269868 330262 270080 330290
rect 270132 330336 270184 330342
rect 270132 330278 270184 330284
rect 269868 161265 269896 330262
rect 270236 316034 270264 330754
rect 269960 316006 270264 316034
rect 269960 161362 269988 316006
rect 269948 161356 270000 161362
rect 269948 161298 270000 161304
rect 269854 161256 269910 161265
rect 269854 161191 269910 161200
rect 269762 160576 269818 160585
rect 269762 160511 269818 160520
rect 269488 158296 269540 158302
rect 269488 158238 269540 158244
rect 269316 155910 269436 155938
rect 269302 155816 269358 155825
rect 269224 155774 269302 155802
rect 269302 155751 269358 155760
rect 269120 155644 269172 155650
rect 269120 155586 269172 155592
rect 268660 155576 268712 155582
rect 268660 155518 268712 155524
rect 265808 155508 265860 155514
rect 265808 155450 265860 155456
rect 260012 155440 260064 155446
rect 260012 155382 260064 155388
rect 260472 155440 260524 155446
rect 269408 155417 269436 155910
rect 270604 155446 270632 337486
rect 270696 333974 270724 337640
rect 271064 337640 271138 337668
rect 271236 337680 271288 337686
rect 270776 337612 270828 337618
rect 270776 337554 270828 337560
rect 270788 336002 270816 337554
rect 270788 335974 271000 336002
rect 270696 333946 270816 333974
rect 270684 330336 270736 330342
rect 270684 330278 270736 330284
rect 270696 155718 270724 330278
rect 270788 155786 270816 333946
rect 270868 330404 270920 330410
rect 270868 330346 270920 330352
rect 270880 155854 270908 330346
rect 270972 158438 271000 335974
rect 271064 330562 271092 337640
rect 271386 337668 271414 338028
rect 271478 337736 271506 338028
rect 271570 337890 271598 338028
rect 271558 337884 271610 337890
rect 271558 337826 271610 337832
rect 271662 337770 271690 338028
rect 271616 337742 271690 337770
rect 271754 337770 271782 338028
rect 271846 337890 271874 338028
rect 271834 337884 271886 337890
rect 271834 337826 271886 337832
rect 271938 337770 271966 338028
rect 271754 337742 271828 337770
rect 271478 337708 271552 337736
rect 271236 337622 271288 337628
rect 271340 337640 271414 337668
rect 271142 337512 271198 337521
rect 271142 337447 271198 337456
rect 271156 330682 271184 337447
rect 271144 330676 271196 330682
rect 271144 330618 271196 330624
rect 271064 330534 271184 330562
rect 271052 330472 271104 330478
rect 271052 330414 271104 330420
rect 270960 158432 271012 158438
rect 270960 158374 271012 158380
rect 271064 158370 271092 330414
rect 271156 158574 271184 330534
rect 271248 161158 271276 337622
rect 271340 330410 271368 337640
rect 271328 330404 271380 330410
rect 271328 330346 271380 330352
rect 271524 325694 271552 337708
rect 271616 330342 271644 337742
rect 271696 337680 271748 337686
rect 271696 337622 271748 337628
rect 271708 336297 271736 337622
rect 271694 336288 271750 336297
rect 271694 336223 271750 336232
rect 271800 335481 271828 337742
rect 271892 337742 271966 337770
rect 271892 337210 271920 337742
rect 272030 337668 272058 338028
rect 272122 337736 272150 338028
rect 272214 337958 272242 338028
rect 272202 337952 272254 337958
rect 272202 337894 272254 337900
rect 272306 337804 272334 338028
rect 272398 337929 272426 338028
rect 272384 337920 272440 337929
rect 272384 337855 272440 337864
rect 272260 337776 272334 337804
rect 272490 337793 272518 338028
rect 272582 337958 272610 338028
rect 272570 337952 272622 337958
rect 272570 337894 272622 337900
rect 272674 337804 272702 338028
rect 272476 337784 272532 337793
rect 272122 337708 272196 337736
rect 272030 337640 272104 337668
rect 271972 337544 272024 337550
rect 271972 337486 272024 337492
rect 271880 337204 271932 337210
rect 271880 337146 271932 337152
rect 271984 337090 272012 337486
rect 271892 337062 272012 337090
rect 271786 335472 271842 335481
rect 271786 335407 271842 335416
rect 271604 330336 271656 330342
rect 271604 330278 271656 330284
rect 271892 325694 271920 337062
rect 271972 333260 272024 333266
rect 271972 333202 272024 333208
rect 271984 328454 272012 333202
rect 272076 331106 272104 337640
rect 272168 333146 272196 337708
rect 272260 333266 272288 337776
rect 272476 337719 272532 337728
rect 272628 337776 272702 337804
rect 272432 337680 272484 337686
rect 272432 337622 272484 337628
rect 272524 337680 272576 337686
rect 272524 337622 272576 337628
rect 272340 337612 272392 337618
rect 272340 337554 272392 337560
rect 272352 335306 272380 337554
rect 272444 336938 272472 337622
rect 272432 336932 272484 336938
rect 272432 336874 272484 336880
rect 272430 336152 272486 336161
rect 272430 336087 272486 336096
rect 272340 335300 272392 335306
rect 272340 335242 272392 335248
rect 272248 333260 272300 333266
rect 272248 333202 272300 333208
rect 272444 333146 272472 336087
rect 272536 333266 272564 337622
rect 272524 333260 272576 333266
rect 272524 333202 272576 333208
rect 272168 333118 272380 333146
rect 272444 333118 272564 333146
rect 272076 331078 272288 331106
rect 272156 331016 272208 331022
rect 272156 330958 272208 330964
rect 271984 328426 272104 328454
rect 271524 325666 271736 325694
rect 271892 325666 272012 325694
rect 271236 161152 271288 161158
rect 271236 161094 271288 161100
rect 271144 158568 271196 158574
rect 271144 158510 271196 158516
rect 271052 158364 271104 158370
rect 271052 158306 271104 158312
rect 270868 155848 270920 155854
rect 270868 155790 270920 155796
rect 270776 155780 270828 155786
rect 270776 155722 270828 155728
rect 270684 155712 270736 155718
rect 270684 155654 270736 155660
rect 271708 155446 271736 325666
rect 271984 158166 272012 325666
rect 272076 158642 272104 328426
rect 272064 158636 272116 158642
rect 272064 158578 272116 158584
rect 272168 158234 272196 330958
rect 272260 158506 272288 331078
rect 272352 161129 272380 333118
rect 272432 333056 272484 333062
rect 272432 332998 272484 333004
rect 272338 161120 272394 161129
rect 272444 161090 272472 332998
rect 272536 161226 272564 333118
rect 272628 333062 272656 337776
rect 272766 337736 272794 338028
rect 272720 337708 272794 337736
rect 272720 335170 272748 337708
rect 272858 337668 272886 338028
rect 272950 337958 272978 338028
rect 272938 337952 272990 337958
rect 272938 337894 272990 337900
rect 273042 337770 273070 338028
rect 273134 337958 273162 338028
rect 273122 337952 273174 337958
rect 273122 337894 273174 337900
rect 273226 337770 273254 338028
rect 273318 337890 273346 338028
rect 273306 337884 273358 337890
rect 273306 337826 273358 337832
rect 273410 337770 273438 338028
rect 273502 337890 273530 338028
rect 273490 337884 273542 337890
rect 273490 337826 273542 337832
rect 273594 337770 273622 338028
rect 273686 337929 273714 338028
rect 273778 337958 273806 338028
rect 273766 337952 273818 337958
rect 273672 337920 273728 337929
rect 273766 337894 273818 337900
rect 273672 337855 273728 337864
rect 273042 337742 273116 337770
rect 273226 337742 273300 337770
rect 272812 337640 272886 337668
rect 272984 337680 273036 337686
rect 272708 335164 272760 335170
rect 272708 335106 272760 335112
rect 272616 333056 272668 333062
rect 272616 332998 272668 333004
rect 272812 331022 272840 337640
rect 272984 337622 273036 337628
rect 272996 332110 273024 337622
rect 272984 332104 273036 332110
rect 272984 332046 273036 332052
rect 272800 331016 272852 331022
rect 272800 330958 272852 330964
rect 273088 325694 273116 337742
rect 273166 337648 273222 337657
rect 273166 337583 273222 337592
rect 273180 335714 273208 337583
rect 273272 336054 273300 337742
rect 273364 337742 273438 337770
rect 273548 337742 273622 337770
rect 273720 337816 273772 337822
rect 273720 337758 273772 337764
rect 273260 336048 273312 336054
rect 273260 335990 273312 335996
rect 273168 335708 273220 335714
rect 273168 335650 273220 335656
rect 273364 326346 273392 337742
rect 273548 333010 273576 337742
rect 273628 337680 273680 337686
rect 273628 337622 273680 337628
rect 273640 336870 273668 337622
rect 273628 336864 273680 336870
rect 273628 336806 273680 336812
rect 273272 326318 273392 326346
rect 273456 332982 273576 333010
rect 273088 325666 273208 325694
rect 272616 163532 272668 163538
rect 272616 163474 272668 163480
rect 272628 162178 272656 163474
rect 272616 162172 272668 162178
rect 272616 162114 272668 162120
rect 272524 161220 272576 161226
rect 272524 161162 272576 161168
rect 272338 161055 272394 161064
rect 272432 161084 272484 161090
rect 272432 161026 272484 161032
rect 272892 158704 272944 158710
rect 272892 158646 272944 158652
rect 272248 158500 272300 158506
rect 272248 158442 272300 158448
rect 272156 158228 272208 158234
rect 272156 158170 272208 158176
rect 271972 158160 272024 158166
rect 271972 158102 272024 158108
rect 272904 155924 272932 158646
rect 271880 155712 271932 155718
rect 271880 155654 271932 155660
rect 271892 155446 271920 155654
rect 270592 155440 270644 155446
rect 260472 155382 260524 155388
rect 269394 155408 269450 155417
rect 270592 155382 270644 155388
rect 271696 155440 271748 155446
rect 271696 155382 271748 155388
rect 271880 155440 271932 155446
rect 273180 155417 273208 325666
rect 273272 156874 273300 326318
rect 273352 325916 273404 325922
rect 273352 325858 273404 325864
rect 273364 163878 273392 325858
rect 273456 163946 273484 332982
rect 273536 332920 273588 332926
rect 273536 332862 273588 332868
rect 273444 163940 273496 163946
rect 273444 163882 273496 163888
rect 273352 163872 273404 163878
rect 273352 163814 273404 163820
rect 273548 163810 273576 332862
rect 273732 328454 273760 337758
rect 273870 337736 273898 338028
rect 273962 337890 273990 338028
rect 274054 337890 274082 338028
rect 274146 337958 274174 338028
rect 274238 337958 274266 338028
rect 274330 337958 274358 338028
rect 274422 337963 274450 338028
rect 274134 337952 274186 337958
rect 274134 337894 274186 337900
rect 274226 337952 274278 337958
rect 274226 337894 274278 337900
rect 274318 337952 274370 337958
rect 274318 337894 274370 337900
rect 274408 337954 274464 337963
rect 274514 337958 274542 338028
rect 273950 337884 274002 337890
rect 273950 337826 274002 337832
rect 274042 337884 274094 337890
rect 274408 337889 274464 337898
rect 274502 337952 274554 337958
rect 274606 337929 274634 338028
rect 274502 337894 274554 337900
rect 274592 337920 274648 337929
rect 274592 337855 274648 337864
rect 274042 337826 274094 337832
rect 274134 337816 274186 337822
rect 274364 337816 274416 337822
rect 274186 337776 274312 337804
rect 274134 337758 274186 337764
rect 273870 337708 273944 337736
rect 273810 337648 273866 337657
rect 273810 337583 273866 337592
rect 273824 334490 273852 337583
rect 273812 334484 273864 334490
rect 273812 334426 273864 334432
rect 273812 333396 273864 333402
rect 273812 333338 273864 333344
rect 273640 328426 273760 328454
rect 273640 174826 273668 328426
rect 273824 326346 273852 333338
rect 273732 326318 273852 326346
rect 273628 174820 273680 174826
rect 273628 174762 273680 174768
rect 273732 174758 273760 326318
rect 273916 325922 273944 337708
rect 274284 337618 274312 337776
rect 274364 337758 274416 337764
rect 274456 337816 274508 337822
rect 274456 337758 274508 337764
rect 274088 337612 274140 337618
rect 274088 337554 274140 337560
rect 274272 337612 274324 337618
rect 274272 337554 274324 337560
rect 273996 337544 274048 337550
rect 273996 337486 274048 337492
rect 273904 325916 273956 325922
rect 273904 325858 273956 325864
rect 274008 325394 274036 337486
rect 274100 332926 274128 337554
rect 274180 337544 274232 337550
rect 274180 337486 274232 337492
rect 274270 337512 274326 337521
rect 274192 333402 274220 337486
rect 274270 337447 274326 337456
rect 274284 335238 274312 337447
rect 274272 335232 274324 335238
rect 274272 335174 274324 335180
rect 274180 333396 274232 333402
rect 274180 333338 274232 333344
rect 274180 333260 274232 333266
rect 274180 333202 274232 333208
rect 274088 332920 274140 332926
rect 274088 332862 274140 332868
rect 274192 328454 274220 333202
rect 274376 333198 274404 337758
rect 274468 333305 274496 337758
rect 274548 337748 274600 337754
rect 274698 337736 274726 338028
rect 274790 337822 274818 338028
rect 274778 337816 274830 337822
rect 274778 337758 274830 337764
rect 274548 337690 274600 337696
rect 274652 337708 274726 337736
rect 274882 337736 274910 338028
rect 274974 337958 275002 338028
rect 274962 337952 275014 337958
rect 274962 337894 275014 337900
rect 275066 337890 275094 338028
rect 275158 337890 275186 338028
rect 275250 337963 275278 338028
rect 275236 337954 275292 337963
rect 275054 337884 275106 337890
rect 275054 337826 275106 337832
rect 275146 337884 275198 337890
rect 275236 337889 275292 337898
rect 275146 337826 275198 337832
rect 275342 337736 275370 338028
rect 275434 337793 275462 338028
rect 275526 337958 275554 338028
rect 275514 337952 275566 337958
rect 275514 337894 275566 337900
rect 275618 337890 275646 338028
rect 275710 337929 275738 338028
rect 275696 337920 275752 337929
rect 275606 337884 275658 337890
rect 275696 337855 275752 337864
rect 275606 337826 275658 337832
rect 275802 337804 275830 338028
rect 275894 337958 275922 338028
rect 275882 337952 275934 337958
rect 275882 337894 275934 337900
rect 275986 337890 276014 338028
rect 275974 337884 276026 337890
rect 275974 337826 276026 337832
rect 274882 337708 274956 337736
rect 274560 334966 274588 337690
rect 274652 337521 274680 337708
rect 274822 337648 274878 337657
rect 274822 337583 274878 337592
rect 274638 337512 274694 337521
rect 274836 337482 274864 337583
rect 274638 337447 274694 337456
rect 274824 337476 274876 337482
rect 274824 337418 274876 337424
rect 274732 337408 274784 337414
rect 274732 337350 274784 337356
rect 274744 336598 274772 337350
rect 274732 336592 274784 336598
rect 274732 336534 274784 336540
rect 274928 335510 274956 337708
rect 275296 337708 275370 337736
rect 275420 337784 275476 337793
rect 275802 337776 275876 337804
rect 275420 337719 275476 337728
rect 275560 337748 275612 337754
rect 275008 337680 275060 337686
rect 275008 337622 275060 337628
rect 274916 335504 274968 335510
rect 274916 335446 274968 335452
rect 275020 335442 275048 337622
rect 275192 337340 275244 337346
rect 275192 337282 275244 337288
rect 275100 337272 275152 337278
rect 275100 337214 275152 337220
rect 274824 335436 274876 335442
rect 274824 335378 274876 335384
rect 275008 335436 275060 335442
rect 275008 335378 275060 335384
rect 274732 335368 274784 335374
rect 274638 335336 274694 335345
rect 274732 335310 274784 335316
rect 274638 335271 274694 335280
rect 274548 334960 274600 334966
rect 274548 334902 274600 334908
rect 274454 333296 274510 333305
rect 274454 333231 274510 333240
rect 274364 333192 274416 333198
rect 274364 333134 274416 333140
rect 273824 325366 274036 325394
rect 274100 328426 274220 328454
rect 273824 179110 273852 325366
rect 274100 321554 274128 328426
rect 274652 328166 274680 335271
rect 274640 328160 274692 328166
rect 274640 328102 274692 328108
rect 274744 326738 274772 335310
rect 274732 326732 274784 326738
rect 274732 326674 274784 326680
rect 274836 326618 274864 335378
rect 275006 335336 275062 335345
rect 275006 335271 275062 335280
rect 273916 321526 274128 321554
rect 274652 326590 274864 326618
rect 273812 179104 273864 179110
rect 273812 179046 273864 179052
rect 273720 174752 273772 174758
rect 273720 174694 273772 174700
rect 273916 169250 273944 321526
rect 273904 169244 273956 169250
rect 273904 169186 273956 169192
rect 273536 163804 273588 163810
rect 273536 163746 273588 163752
rect 274652 163674 274680 326590
rect 274732 326460 274784 326466
rect 274732 326402 274784 326408
rect 274744 165306 274772 326402
rect 275020 326346 275048 335271
rect 274836 326318 275048 326346
rect 274732 165300 274784 165306
rect 274732 165242 274784 165248
rect 274836 165238 274864 326318
rect 274916 326188 274968 326194
rect 274916 326130 274968 326136
rect 274824 165232 274876 165238
rect 274824 165174 274876 165180
rect 274928 165170 274956 326130
rect 275008 326120 275060 326126
rect 275008 326062 275060 326068
rect 274916 165164 274968 165170
rect 274916 165106 274968 165112
rect 275020 165102 275048 326062
rect 275112 174690 275140 337214
rect 275204 326482 275232 337282
rect 275296 326602 275324 337708
rect 275848 337736 275876 337776
rect 276078 337770 276106 338028
rect 276170 337958 276198 338028
rect 276262 337958 276290 338028
rect 276354 337958 276382 338028
rect 276158 337952 276210 337958
rect 276158 337894 276210 337900
rect 276250 337952 276302 337958
rect 276250 337894 276302 337900
rect 276342 337952 276394 337958
rect 276342 337894 276394 337900
rect 276204 337816 276256 337822
rect 276078 337742 276152 337770
rect 276446 337793 276474 338028
rect 276538 337958 276566 338028
rect 276630 337958 276658 338028
rect 276526 337952 276578 337958
rect 276526 337894 276578 337900
rect 276618 337952 276670 337958
rect 276618 337894 276670 337900
rect 276204 337758 276256 337764
rect 276432 337784 276488 337793
rect 275848 337708 275968 337736
rect 275560 337690 275612 337696
rect 275468 337680 275520 337686
rect 275468 337622 275520 337628
rect 275376 337612 275428 337618
rect 275376 337554 275428 337560
rect 275388 335374 275416 337554
rect 275376 335368 275428 335374
rect 275376 335310 275428 335316
rect 275284 326596 275336 326602
rect 275284 326538 275336 326544
rect 275204 326454 275416 326482
rect 275192 326392 275244 326398
rect 275192 326334 275244 326340
rect 275204 176390 275232 326334
rect 275284 326256 275336 326262
rect 275284 326198 275336 326204
rect 275192 176384 275244 176390
rect 275192 176326 275244 176332
rect 275296 176322 275324 326198
rect 275388 176458 275416 326454
rect 275480 326194 275508 337622
rect 275572 326262 275600 337690
rect 275744 337680 275796 337686
rect 275744 337622 275796 337628
rect 275834 337648 275890 337657
rect 275650 337512 275706 337521
rect 275650 337447 275706 337456
rect 275664 330614 275692 337447
rect 275756 337142 275784 337622
rect 275834 337583 275890 337592
rect 275744 337136 275796 337142
rect 275744 337078 275796 337084
rect 275848 335374 275876 337583
rect 275836 335368 275888 335374
rect 275836 335310 275888 335316
rect 275940 332594 275968 337708
rect 276020 337612 276072 337618
rect 276020 337554 276072 337560
rect 276032 336394 276060 337554
rect 276124 337006 276152 337742
rect 276112 337000 276164 337006
rect 276112 336942 276164 336948
rect 276020 336388 276072 336394
rect 276020 336330 276072 336336
rect 276216 335578 276244 337758
rect 276722 337770 276750 338028
rect 276814 337958 276842 338028
rect 276906 337958 276934 338028
rect 276998 337958 277026 338028
rect 277090 337963 277118 338028
rect 276802 337952 276854 337958
rect 276802 337894 276854 337900
rect 276894 337952 276946 337958
rect 276894 337894 276946 337900
rect 276986 337952 277038 337958
rect 276986 337894 277038 337900
rect 277076 337954 277132 337963
rect 277076 337889 277132 337898
rect 276848 337816 276900 337822
rect 276722 337742 276796 337770
rect 276848 337758 276900 337764
rect 276432 337719 276488 337728
rect 276296 337680 276348 337686
rect 276664 337680 276716 337686
rect 276296 337622 276348 337628
rect 276478 337648 276534 337657
rect 276204 335572 276256 335578
rect 276204 335514 276256 335520
rect 276112 335436 276164 335442
rect 276112 335378 276164 335384
rect 275848 332566 275968 332594
rect 275652 330608 275704 330614
rect 275652 330550 275704 330556
rect 275652 328160 275704 328166
rect 275652 328102 275704 328108
rect 275560 326256 275612 326262
rect 275560 326198 275612 326204
rect 275468 326188 275520 326194
rect 275468 326130 275520 326136
rect 275664 325038 275692 328102
rect 275848 326126 275876 332566
rect 276020 326392 276072 326398
rect 276020 326334 276072 326340
rect 275836 326120 275888 326126
rect 275836 326062 275888 326068
rect 275652 325032 275704 325038
rect 275652 324974 275704 324980
rect 275376 176452 275428 176458
rect 275376 176394 275428 176400
rect 275284 176316 275336 176322
rect 275284 176258 275336 176264
rect 275100 174684 275152 174690
rect 275100 174626 275152 174632
rect 275008 165096 275060 165102
rect 275008 165038 275060 165044
rect 276032 164898 276060 326334
rect 276124 164966 276152 335378
rect 276308 327418 276336 337622
rect 276664 337622 276716 337628
rect 276478 337583 276534 337592
rect 276388 337476 276440 337482
rect 276388 337418 276440 337424
rect 276296 327412 276348 327418
rect 276296 327354 276348 327360
rect 276400 326346 276428 337418
rect 276492 333538 276520 337583
rect 276572 337544 276624 337550
rect 276572 337486 276624 337492
rect 276584 333713 276612 337486
rect 276676 335442 276704 337622
rect 276664 335436 276716 335442
rect 276664 335378 276716 335384
rect 276768 335322 276796 337742
rect 276676 335294 276796 335322
rect 276570 333704 276626 333713
rect 276570 333639 276626 333648
rect 276480 333532 276532 333538
rect 276480 333474 276532 333480
rect 276572 333192 276624 333198
rect 276572 333134 276624 333140
rect 276584 326346 276612 333134
rect 276216 326318 276428 326346
rect 276492 326318 276612 326346
rect 276216 165034 276244 326318
rect 276296 326256 276348 326262
rect 276296 326198 276348 326204
rect 276308 176254 276336 326198
rect 276492 321554 276520 326318
rect 276676 326262 276704 335294
rect 276756 334484 276808 334490
rect 276756 334426 276808 334432
rect 276664 326256 276716 326262
rect 276664 326198 276716 326204
rect 276492 321526 276704 321554
rect 276296 176248 276348 176254
rect 276296 176190 276348 176196
rect 276204 165028 276256 165034
rect 276204 164970 276256 164976
rect 276112 164960 276164 164966
rect 276112 164902 276164 164908
rect 276020 164892 276072 164898
rect 276020 164834 276072 164840
rect 274640 163668 274692 163674
rect 274640 163610 274692 163616
rect 276676 162314 276704 321526
rect 276768 170814 276796 334426
rect 276860 326398 276888 337758
rect 276940 337748 276992 337754
rect 276940 337690 276992 337696
rect 276952 333470 276980 337690
rect 277032 337680 277084 337686
rect 277182 337668 277210 338028
rect 277274 337958 277302 338028
rect 277262 337952 277314 337958
rect 277262 337894 277314 337900
rect 277366 337736 277394 338028
rect 277320 337708 277394 337736
rect 277458 337736 277486 338028
rect 277550 337804 277578 338028
rect 277642 337958 277670 338028
rect 277630 337952 277682 337958
rect 277630 337894 277682 337900
rect 277734 337804 277762 338028
rect 277826 337958 277854 338028
rect 277918 337958 277946 338028
rect 278010 337958 278038 338028
rect 278102 337958 278130 338028
rect 278194 337958 278222 338028
rect 278286 337963 278314 338028
rect 277814 337952 277866 337958
rect 277814 337894 277866 337900
rect 277906 337952 277958 337958
rect 277906 337894 277958 337900
rect 277998 337952 278050 337958
rect 277998 337894 278050 337900
rect 278090 337952 278142 337958
rect 278090 337894 278142 337900
rect 278182 337952 278234 337958
rect 278182 337894 278234 337900
rect 278272 337954 278328 337963
rect 278272 337889 278328 337898
rect 278378 337822 278406 338028
rect 278044 337816 278096 337822
rect 277550 337776 277624 337804
rect 277734 337776 277808 337804
rect 277458 337708 277532 337736
rect 277182 337640 277256 337668
rect 277032 337622 277084 337628
rect 276940 333464 276992 333470
rect 276940 333406 276992 333412
rect 277044 328454 277072 337622
rect 277124 337544 277176 337550
rect 277124 337486 277176 337492
rect 277136 336025 277164 337486
rect 277228 336938 277256 337640
rect 277216 336932 277268 336938
rect 277216 336874 277268 336880
rect 277320 336784 277348 337708
rect 277320 336756 277440 336784
rect 277308 336660 277360 336666
rect 277308 336602 277360 336608
rect 277122 336016 277178 336025
rect 277122 335951 277178 335960
rect 277320 335646 277348 336602
rect 277412 336462 277440 336756
rect 277400 336456 277452 336462
rect 277400 336398 277452 336404
rect 277400 335912 277452 335918
rect 277400 335854 277452 335860
rect 277308 335640 277360 335646
rect 277308 335582 277360 335588
rect 276952 328426 277072 328454
rect 276952 327894 276980 328426
rect 276940 327888 276992 327894
rect 276940 327830 276992 327836
rect 276940 327412 276992 327418
rect 276940 327354 276992 327360
rect 276848 326392 276900 326398
rect 276848 326334 276900 326340
rect 276952 323610 276980 327354
rect 276940 323604 276992 323610
rect 276940 323546 276992 323552
rect 276756 170808 276808 170814
rect 276756 170750 276808 170756
rect 277412 166530 277440 335854
rect 277504 326346 277532 337708
rect 277596 336190 277624 337776
rect 277676 337680 277728 337686
rect 277676 337622 277728 337628
rect 277584 336184 277636 336190
rect 277584 336126 277636 336132
rect 277584 333260 277636 333266
rect 277584 333202 277636 333208
rect 277596 326466 277624 333202
rect 277688 326466 277716 337622
rect 277780 335918 277808 337776
rect 278366 337816 278418 337822
rect 278044 337758 278096 337764
rect 278226 337784 278282 337793
rect 277952 337612 278004 337618
rect 277952 337554 278004 337560
rect 277860 337544 277912 337550
rect 277860 337486 277912 337492
rect 277768 335912 277820 335918
rect 277768 335854 277820 335860
rect 277872 333974 277900 337486
rect 277780 333946 277900 333974
rect 277584 326460 277636 326466
rect 277584 326402 277636 326408
rect 277676 326460 277728 326466
rect 277676 326402 277728 326408
rect 277780 326346 277808 333946
rect 277860 326460 277912 326466
rect 277860 326402 277912 326408
rect 277504 326318 277624 326346
rect 277492 326188 277544 326194
rect 277492 326130 277544 326136
rect 277400 166524 277452 166530
rect 277400 166466 277452 166472
rect 277504 166462 277532 326130
rect 277596 166666 277624 326318
rect 277688 326318 277808 326346
rect 277688 176186 277716 326318
rect 277768 326256 277820 326262
rect 277768 326198 277820 326204
rect 277676 176180 277728 176186
rect 277676 176122 277728 176128
rect 277780 176050 277808 326198
rect 277872 178974 277900 326402
rect 277964 180198 277992 337554
rect 278056 333974 278084 337758
rect 278366 337758 278418 337764
rect 278226 337719 278282 337728
rect 278470 337736 278498 338028
rect 278562 337963 278590 338028
rect 278548 337954 278604 337963
rect 278548 337889 278604 337898
rect 278654 337793 278682 338028
rect 278746 337958 278774 338028
rect 278734 337952 278786 337958
rect 278838 337929 278866 338028
rect 278930 337958 278958 338028
rect 279022 337958 279050 338028
rect 279114 337958 279142 338028
rect 279206 337958 279234 338028
rect 279298 337958 279326 338028
rect 278918 337952 278970 337958
rect 278734 337894 278786 337900
rect 278824 337920 278880 337929
rect 278918 337894 278970 337900
rect 279010 337952 279062 337958
rect 279010 337894 279062 337900
rect 279102 337952 279154 337958
rect 279102 337894 279154 337900
rect 279194 337952 279246 337958
rect 279194 337894 279246 337900
rect 279286 337952 279338 337958
rect 279286 337894 279338 337900
rect 278824 337855 278880 337864
rect 278780 337816 278832 337822
rect 278640 337784 278696 337793
rect 278136 337476 278188 337482
rect 278136 337418 278188 337424
rect 278148 335986 278176 337418
rect 278136 335980 278188 335986
rect 278136 335922 278188 335928
rect 278056 333946 278176 333974
rect 278148 326194 278176 333946
rect 278240 327826 278268 337719
rect 278470 337708 278544 337736
rect 278780 337758 278832 337764
rect 278640 337719 278696 337728
rect 278320 337680 278372 337686
rect 278320 337622 278372 337628
rect 278410 337648 278466 337657
rect 278332 333266 278360 337622
rect 278410 337583 278466 337592
rect 278424 333577 278452 337583
rect 278410 333568 278466 333577
rect 278410 333503 278466 333512
rect 278516 333305 278544 337708
rect 278596 337680 278648 337686
rect 278596 337622 278648 337628
rect 278688 337680 278740 337686
rect 278688 337622 278740 337628
rect 278608 335918 278636 337622
rect 278700 336530 278728 337622
rect 278688 336524 278740 336530
rect 278688 336466 278740 336472
rect 278596 335912 278648 335918
rect 278596 335854 278648 335860
rect 278502 333296 278558 333305
rect 278320 333260 278372 333266
rect 278502 333231 278558 333240
rect 278320 333202 278372 333208
rect 278228 327820 278280 327826
rect 278228 327762 278280 327768
rect 278136 326188 278188 326194
rect 278136 326130 278188 326136
rect 278792 325582 278820 337758
rect 278964 337748 279016 337754
rect 279390 337736 279418 338028
rect 279482 337958 279510 338028
rect 279574 337958 279602 338028
rect 279666 337958 279694 338028
rect 279470 337952 279522 337958
rect 279470 337894 279522 337900
rect 279562 337952 279614 337958
rect 279562 337894 279614 337900
rect 279654 337952 279706 337958
rect 279654 337894 279706 337900
rect 279516 337748 279568 337754
rect 279390 337708 279464 337736
rect 278964 337690 279016 337696
rect 278872 337612 278924 337618
rect 278872 337554 278924 337560
rect 278780 325576 278832 325582
rect 278780 325518 278832 325524
rect 278780 325440 278832 325446
rect 278780 325382 278832 325388
rect 277952 180192 278004 180198
rect 277952 180134 278004 180140
rect 277860 178968 277912 178974
rect 277860 178910 277912 178916
rect 277768 176044 277820 176050
rect 277768 175986 277820 175992
rect 277584 166660 277636 166666
rect 277584 166602 277636 166608
rect 277492 166456 277544 166462
rect 277492 166398 277544 166404
rect 278792 166394 278820 325382
rect 278884 168162 278912 337554
rect 278976 336274 279004 337690
rect 279240 337612 279292 337618
rect 279240 337554 279292 337560
rect 279332 337612 279384 337618
rect 279332 337554 279384 337560
rect 279148 337544 279200 337550
rect 279148 337486 279200 337492
rect 278976 336246 279096 336274
rect 278964 336184 279016 336190
rect 278964 336126 279016 336132
rect 278976 333402 279004 336126
rect 278964 333396 279016 333402
rect 278964 333338 279016 333344
rect 279068 328454 279096 336246
rect 279160 333334 279188 337486
rect 279148 333328 279200 333334
rect 279148 333270 279200 333276
rect 279068 328426 279188 328454
rect 278964 326392 279016 326398
rect 278964 326334 279016 326340
rect 278872 168156 278924 168162
rect 278872 168098 278924 168104
rect 278976 168026 279004 326334
rect 279056 325848 279108 325854
rect 279056 325790 279108 325796
rect 279068 168094 279096 325790
rect 279160 170678 279188 328426
rect 279148 170672 279200 170678
rect 279148 170614 279200 170620
rect 279252 170610 279280 337554
rect 279344 335850 279372 337554
rect 279332 335844 279384 335850
rect 279332 335786 279384 335792
rect 279436 333974 279464 337708
rect 279516 337690 279568 337696
rect 279608 337748 279660 337754
rect 279758 337736 279786 338028
rect 279850 337958 279878 338028
rect 279838 337952 279890 337958
rect 279942 337929 279970 338028
rect 280034 337958 280062 338028
rect 280022 337952 280074 337958
rect 279838 337894 279890 337900
rect 279928 337920 279984 337929
rect 280022 337894 280074 337900
rect 280126 337895 280154 338028
rect 280218 337958 280246 338028
rect 280206 337952 280258 337958
rect 279928 337855 279984 337864
rect 280112 337886 280168 337895
rect 280206 337894 280258 337900
rect 279976 337816 280028 337822
rect 280112 337821 280168 337830
rect 279608 337690 279660 337696
rect 279712 337708 279786 337736
rect 279974 337784 279976 337793
rect 280028 337784 280030 337793
rect 280310 337736 280338 338028
rect 280402 337929 280430 338028
rect 280388 337920 280444 337929
rect 280494 337890 280522 338028
rect 280586 337890 280614 338028
rect 280388 337855 280444 337864
rect 280482 337884 280534 337890
rect 280482 337826 280534 337832
rect 280574 337884 280626 337890
rect 280574 337826 280626 337832
rect 280678 337770 280706 338028
rect 280770 337804 280798 338028
rect 280862 337963 280890 338028
rect 280848 337954 280904 337963
rect 280848 337889 280904 337898
rect 280954 337890 280982 338028
rect 281046 337958 281074 338028
rect 281034 337952 281086 337958
rect 281034 337894 281086 337900
rect 281138 337890 281166 338028
rect 280942 337884 280994 337890
rect 280942 337826 280994 337832
rect 281126 337884 281178 337890
rect 281126 337826 281178 337832
rect 281230 337822 281258 338028
rect 281322 337890 281350 338028
rect 281414 337958 281442 338028
rect 281402 337952 281454 337958
rect 281506 337929 281534 338028
rect 281402 337894 281454 337900
rect 281492 337920 281548 337929
rect 281310 337884 281362 337890
rect 281598 337890 281626 338028
rect 281492 337855 281548 337864
rect 281586 337884 281638 337890
rect 281310 337826 281362 337832
rect 281586 337826 281638 337832
rect 281218 337816 281270 337822
rect 280770 337776 280844 337804
rect 279974 337719 280030 337728
rect 280264 337708 280338 337736
rect 280632 337742 280706 337770
rect 279344 333946 279464 333974
rect 279344 325854 279372 333946
rect 279332 325848 279384 325854
rect 279332 325790 279384 325796
rect 279528 325786 279556 337690
rect 279620 326398 279648 337690
rect 279608 326392 279660 326398
rect 279608 326334 279660 326340
rect 279516 325780 279568 325786
rect 279516 325722 279568 325728
rect 279712 325666 279740 337708
rect 279792 337544 279844 337550
rect 279792 337486 279844 337492
rect 279804 336598 279832 337486
rect 279884 337476 279936 337482
rect 279884 337418 279936 337424
rect 279792 336592 279844 336598
rect 279792 336534 279844 336540
rect 279896 336410 279924 337418
rect 280068 337408 280120 337414
rect 280068 337350 280120 337356
rect 279804 336382 279924 336410
rect 279804 333441 279832 336382
rect 279882 336288 279938 336297
rect 279882 336223 279884 336232
rect 279936 336223 279938 336232
rect 279884 336194 279936 336200
rect 279884 334960 279936 334966
rect 279884 334902 279936 334908
rect 279790 333432 279846 333441
rect 279790 333367 279846 333376
rect 279896 326670 279924 334902
rect 280080 333266 280108 337350
rect 280264 337278 280292 337708
rect 280528 337680 280580 337686
rect 280528 337622 280580 337628
rect 280344 337612 280396 337618
rect 280344 337554 280396 337560
rect 280436 337612 280488 337618
rect 280436 337554 280488 337560
rect 280252 337272 280304 337278
rect 280252 337214 280304 337220
rect 280356 336870 280384 337554
rect 280344 336864 280396 336870
rect 280344 336806 280396 336812
rect 280252 336796 280304 336802
rect 280252 336738 280304 336744
rect 280068 333260 280120 333266
rect 280068 333202 280120 333208
rect 279884 326664 279936 326670
rect 279884 326606 279936 326612
rect 279344 325638 279740 325666
rect 279240 170604 279292 170610
rect 279240 170546 279292 170552
rect 279344 170542 279372 325638
rect 279424 325576 279476 325582
rect 279424 325518 279476 325524
rect 279436 175982 279464 325518
rect 279424 175976 279476 175982
rect 279424 175918 279476 175924
rect 279332 170536 279384 170542
rect 279332 170478 279384 170484
rect 279056 168088 279108 168094
rect 279056 168030 279108 168036
rect 278964 168020 279016 168026
rect 278964 167962 279016 167968
rect 280264 167822 280292 336738
rect 280342 336696 280398 336705
rect 280342 336631 280398 336640
rect 280356 167958 280384 336631
rect 280344 167952 280396 167958
rect 280344 167894 280396 167900
rect 280448 167890 280476 337554
rect 280540 326482 280568 337622
rect 280632 326618 280660 337742
rect 280816 337600 280844 337776
rect 281690 337770 281718 338028
rect 281782 337958 281810 338028
rect 281770 337952 281822 337958
rect 281770 337894 281822 337900
rect 281218 337758 281270 337764
rect 281080 337748 281132 337754
rect 281080 337690 281132 337696
rect 281460 337742 281718 337770
rect 280988 337612 281040 337618
rect 280816 337572 280936 337600
rect 280804 337476 280856 337482
rect 280804 337418 280856 337424
rect 280712 336320 280764 336326
rect 280710 336288 280712 336297
rect 280764 336288 280766 336297
rect 280710 336223 280766 336232
rect 280816 333305 280844 337418
rect 280908 336841 280936 337572
rect 280988 337554 281040 337560
rect 280894 336832 280950 336841
rect 280894 336767 280950 336776
rect 280894 336696 280950 336705
rect 280894 336631 280950 336640
rect 280802 333296 280858 333305
rect 280802 333231 280858 333240
rect 280632 326590 280844 326618
rect 280540 326454 280752 326482
rect 280528 326392 280580 326398
rect 280528 326334 280580 326340
rect 280540 169182 280568 326334
rect 280620 326324 280672 326330
rect 280620 326266 280672 326272
rect 280632 174622 280660 326266
rect 280724 177818 280752 326454
rect 280816 326330 280844 326590
rect 280804 326324 280856 326330
rect 280804 326266 280856 326272
rect 280908 324970 280936 336631
rect 281000 335753 281028 337554
rect 280986 335744 281042 335753
rect 280986 335679 281042 335688
rect 280896 324964 280948 324970
rect 280896 324906 280948 324912
rect 281092 321554 281120 337690
rect 281354 337648 281410 337657
rect 281172 337612 281224 337618
rect 281354 337583 281410 337592
rect 281172 337554 281224 337560
rect 281184 336802 281212 337554
rect 281264 337544 281316 337550
rect 281264 337486 281316 337492
rect 281172 336796 281224 336802
rect 281172 336738 281224 336744
rect 281276 326398 281304 337486
rect 281368 336190 281396 337583
rect 281460 337414 281488 337742
rect 281874 337736 281902 338028
rect 281966 337890 281994 338028
rect 282058 337929 282086 338028
rect 282150 337958 282178 338028
rect 282242 337958 282270 338028
rect 282138 337952 282190 337958
rect 282044 337920 282100 337929
rect 281954 337884 282006 337890
rect 282138 337894 282190 337900
rect 282230 337952 282282 337958
rect 282334 337929 282362 338028
rect 282230 337894 282282 337900
rect 282320 337920 282376 337929
rect 282044 337855 282100 337864
rect 282320 337855 282376 337864
rect 281954 337826 282006 337832
rect 281828 337708 281902 337736
rect 281998 337784 282054 337793
rect 281998 337719 282054 337728
rect 282092 337748 282144 337754
rect 281540 337680 281592 337686
rect 281540 337622 281592 337628
rect 281448 337408 281500 337414
rect 281448 337350 281500 337356
rect 281448 337272 281500 337278
rect 281448 337214 281500 337220
rect 281356 336184 281408 336190
rect 281356 336126 281408 336132
rect 281356 335640 281408 335646
rect 281356 335582 281408 335588
rect 281368 330682 281396 335582
rect 281356 330676 281408 330682
rect 281356 330618 281408 330624
rect 281264 326392 281316 326398
rect 281264 326334 281316 326340
rect 280816 321526 281120 321554
rect 280712 177812 280764 177818
rect 280712 177754 280764 177760
rect 280816 177750 280844 321526
rect 280804 177744 280856 177750
rect 280804 177686 280856 177692
rect 280620 174616 280672 174622
rect 280620 174558 280672 174564
rect 280528 169176 280580 169182
rect 280528 169118 280580 169124
rect 280436 167884 280488 167890
rect 280436 167826 280488 167832
rect 280252 167816 280304 167822
rect 280252 167758 280304 167764
rect 278780 166388 278832 166394
rect 278780 166330 278832 166336
rect 276664 162308 276716 162314
rect 276664 162250 276716 162256
rect 281460 161022 281488 337214
rect 281552 336258 281580 337622
rect 281632 337612 281684 337618
rect 281632 337554 281684 337560
rect 281540 336252 281592 336258
rect 281540 336194 281592 336200
rect 281540 336116 281592 336122
rect 281540 336058 281592 336064
rect 281448 161016 281500 161022
rect 281448 160958 281500 160964
rect 277398 158400 277454 158409
rect 277398 158335 277454 158344
rect 273260 156868 273312 156874
rect 273260 156810 273312 156816
rect 277412 155924 277440 158335
rect 281264 158024 281316 158030
rect 281264 157966 281316 157972
rect 281276 155924 281304 157966
rect 281552 156806 281580 336058
rect 281644 159526 281672 337554
rect 281724 336796 281776 336802
rect 281724 336738 281776 336744
rect 281736 160954 281764 336738
rect 281828 336002 281856 337708
rect 281908 337272 281960 337278
rect 281908 337214 281960 337220
rect 281920 336841 281948 337214
rect 281906 336832 281962 336841
rect 281906 336767 281962 336776
rect 281828 335974 281948 336002
rect 281816 335504 281868 335510
rect 281816 335446 281868 335452
rect 281828 332042 281856 335446
rect 281816 332036 281868 332042
rect 281816 331978 281868 331984
rect 281816 322652 281868 322658
rect 281816 322594 281868 322600
rect 281828 167754 281856 322594
rect 281920 169114 281948 335974
rect 282012 326466 282040 337719
rect 282426 337736 282454 338028
rect 282092 337690 282144 337696
rect 282380 337708 282454 337736
rect 282518 337736 282546 338028
rect 282610 337890 282638 338028
rect 282598 337884 282650 337890
rect 282598 337826 282650 337832
rect 282702 337736 282730 338028
rect 282794 337929 282822 338028
rect 282780 337920 282836 337929
rect 282886 337890 282914 338028
rect 282978 337958 283006 338028
rect 282966 337952 283018 337958
rect 282966 337894 283018 337900
rect 282780 337855 282836 337864
rect 282874 337884 282926 337890
rect 282874 337826 282926 337832
rect 283070 337770 283098 338028
rect 283162 337822 283190 338028
rect 283024 337742 283098 337770
rect 283150 337816 283202 337822
rect 283150 337758 283202 337764
rect 282518 337708 282592 337736
rect 282702 337708 282776 337736
rect 282000 326460 282052 326466
rect 282000 326402 282052 326408
rect 282104 326346 282132 337690
rect 282276 337680 282328 337686
rect 282276 337622 282328 337628
rect 282288 336122 282316 337622
rect 282276 336116 282328 336122
rect 282276 336058 282328 336064
rect 282380 331214 282408 337708
rect 282460 337340 282512 337346
rect 282460 337282 282512 337288
rect 282472 333849 282500 337282
rect 282564 336802 282592 337708
rect 282644 337612 282696 337618
rect 282644 337554 282696 337560
rect 282552 336796 282604 336802
rect 282552 336738 282604 336744
rect 282656 335354 282684 337554
rect 282748 336297 282776 337708
rect 282918 337512 282974 337521
rect 282918 337447 282974 337456
rect 282734 336288 282790 336297
rect 282734 336223 282790 336232
rect 282564 335326 282684 335354
rect 282458 333840 282514 333849
rect 282458 333775 282514 333784
rect 282012 326318 282132 326346
rect 282196 331186 282408 331214
rect 282012 170474 282040 326318
rect 282196 326210 282224 331186
rect 282276 326460 282328 326466
rect 282276 326402 282328 326408
rect 282104 326182 282224 326210
rect 282000 170468 282052 170474
rect 282000 170410 282052 170416
rect 282104 170406 282132 326182
rect 282288 321554 282316 326402
rect 282564 322658 282592 335326
rect 282552 322652 282604 322658
rect 282552 322594 282604 322600
rect 282196 321526 282316 321554
rect 282932 321554 282960 337447
rect 283024 328438 283052 337742
rect 283104 337680 283156 337686
rect 283254 337668 283282 338028
rect 283346 337890 283374 338028
rect 283334 337884 283386 337890
rect 283334 337826 283386 337832
rect 283438 337770 283466 338028
rect 283104 337622 283156 337628
rect 283208 337640 283282 337668
rect 283392 337742 283466 337770
rect 283012 328432 283064 328438
rect 283012 328374 283064 328380
rect 282932 321526 283052 321554
rect 282196 184210 282224 321526
rect 282184 184204 282236 184210
rect 282184 184146 282236 184152
rect 282092 170400 282144 170406
rect 282092 170342 282144 170348
rect 281908 169108 281960 169114
rect 281908 169050 281960 169056
rect 281816 167748 281868 167754
rect 281816 167690 281868 167696
rect 281724 160948 281776 160954
rect 281724 160890 281776 160896
rect 281632 159520 281684 159526
rect 281632 159462 281684 159468
rect 281540 156800 281592 156806
rect 281540 156742 281592 156748
rect 283024 156738 283052 321526
rect 283116 169046 283144 337622
rect 283208 336705 283236 337640
rect 283288 337544 283340 337550
rect 283288 337486 283340 337492
rect 283194 336696 283250 336705
rect 283194 336631 283250 336640
rect 283196 336184 283248 336190
rect 283196 336126 283248 336132
rect 283208 335782 283236 336126
rect 283196 335776 283248 335782
rect 283196 335718 283248 335724
rect 283196 334620 283248 334626
rect 283196 334562 283248 334568
rect 283208 172038 283236 334562
rect 283300 172106 283328 337486
rect 283392 334626 283420 337742
rect 283530 337736 283558 338028
rect 283622 337890 283650 338028
rect 283610 337884 283662 337890
rect 283610 337826 283662 337832
rect 283530 337708 283604 337736
rect 283472 337544 283524 337550
rect 283472 337486 283524 337492
rect 283484 336841 283512 337486
rect 283576 337464 283604 337708
rect 283714 337668 283742 338028
rect 283806 337736 283834 338028
rect 283898 337929 283926 338028
rect 283990 337958 284018 338028
rect 283978 337952 284030 337958
rect 283884 337920 283940 337929
rect 283978 337894 284030 337900
rect 283884 337855 283940 337864
rect 284082 337822 284110 338028
rect 283932 337816 283984 337822
rect 283932 337758 283984 337764
rect 284070 337816 284122 337822
rect 284070 337758 284122 337764
rect 283806 337708 283880 337736
rect 283714 337640 283788 337668
rect 283576 337436 283696 337464
rect 283564 337340 283616 337346
rect 283564 337282 283616 337288
rect 283470 336832 283526 336841
rect 283470 336767 283526 336776
rect 283470 335472 283526 335481
rect 283470 335407 283526 335416
rect 283484 335102 283512 335407
rect 283472 335096 283524 335102
rect 283472 335038 283524 335044
rect 283380 334620 283432 334626
rect 283380 334562 283432 334568
rect 283576 331214 283604 337282
rect 283392 331186 283604 331214
rect 283288 172100 283340 172106
rect 283288 172042 283340 172048
rect 283196 172032 283248 172038
rect 283196 171974 283248 171980
rect 283392 171970 283420 331186
rect 283668 329186 283696 337436
rect 283760 337414 283788 337640
rect 283748 337408 283800 337414
rect 283748 337350 283800 337356
rect 283748 337272 283800 337278
rect 283748 337214 283800 337220
rect 283760 336190 283788 337214
rect 283748 336184 283800 336190
rect 283748 336126 283800 336132
rect 283748 335368 283800 335374
rect 283748 335310 283800 335316
rect 283656 329180 283708 329186
rect 283656 329122 283708 329128
rect 283472 328432 283524 328438
rect 283472 328374 283524 328380
rect 283484 172174 283512 328374
rect 283760 316034 283788 335310
rect 283852 331214 283880 337708
rect 283944 335481 283972 337758
rect 284024 337680 284076 337686
rect 284174 337668 284202 338028
rect 284266 337822 284294 338028
rect 284358 337958 284386 338028
rect 284346 337952 284398 337958
rect 284450 337929 284478 338028
rect 284542 337958 284570 338028
rect 284530 337952 284582 337958
rect 284346 337894 284398 337900
rect 284436 337920 284492 337929
rect 284530 337894 284582 337900
rect 284634 337890 284662 338028
rect 284726 337890 284754 338028
rect 284436 337855 284492 337864
rect 284622 337884 284674 337890
rect 284622 337826 284674 337832
rect 284714 337884 284766 337890
rect 284714 337826 284766 337832
rect 284254 337816 284306 337822
rect 284254 337758 284306 337764
rect 284484 337748 284536 337754
rect 284818 337736 284846 338028
rect 284484 337690 284536 337696
rect 284772 337708 284846 337736
rect 284024 337622 284076 337628
rect 284128 337640 284202 337668
rect 284298 337648 284354 337657
rect 284036 335889 284064 337622
rect 284022 335880 284078 335889
rect 284022 335815 284078 335824
rect 284128 335481 284156 337640
rect 284298 337583 284354 337592
rect 284392 337612 284444 337618
rect 284208 337544 284260 337550
rect 284208 337486 284260 337492
rect 284220 335617 284248 337486
rect 284206 335608 284262 335617
rect 284206 335543 284262 335552
rect 283930 335472 283986 335481
rect 283930 335407 283986 335416
rect 284114 335472 284170 335481
rect 284114 335407 284170 335416
rect 283852 331186 284064 331214
rect 283576 316006 283788 316034
rect 283576 179042 283604 316006
rect 283564 179036 283616 179042
rect 283564 178978 283616 178984
rect 283472 172168 283524 172174
rect 283472 172110 283524 172116
rect 283380 171964 283432 171970
rect 283380 171906 283432 171912
rect 283104 169040 283156 169046
rect 283104 168982 283156 168988
rect 283012 156732 283064 156738
rect 283012 156674 283064 156680
rect 284036 155689 284064 331186
rect 284312 326738 284340 337583
rect 284392 337554 284444 337560
rect 284404 336122 284432 337554
rect 284392 336116 284444 336122
rect 284392 336058 284444 336064
rect 284392 334620 284444 334626
rect 284392 334562 284444 334568
rect 284300 326732 284352 326738
rect 284300 326674 284352 326680
rect 284404 158001 284432 334562
rect 284496 326466 284524 337690
rect 284576 337680 284628 337686
rect 284576 337622 284628 337628
rect 284484 326460 284536 326466
rect 284484 326402 284536 326408
rect 284588 326346 284616 337622
rect 284668 337612 284720 337618
rect 284668 337554 284720 337560
rect 284496 326318 284616 326346
rect 284496 158098 284524 326318
rect 284576 326256 284628 326262
rect 284576 326198 284628 326204
rect 284588 162246 284616 326198
rect 284680 171902 284708 337554
rect 284772 326262 284800 337708
rect 284910 337668 284938 338028
rect 285002 337793 285030 338028
rect 284988 337784 285044 337793
rect 284988 337719 285044 337728
rect 284864 337640 284938 337668
rect 284864 334626 284892 337640
rect 285094 337634 285122 338028
rect 285186 337890 285214 338028
rect 285278 337958 285306 338028
rect 285266 337952 285318 337958
rect 285266 337894 285318 337900
rect 285370 337890 285398 338028
rect 285462 337890 285490 338028
rect 285554 337890 285582 338028
rect 285646 337929 285674 338028
rect 285632 337920 285688 337929
rect 285174 337884 285226 337890
rect 285174 337826 285226 337832
rect 285358 337884 285410 337890
rect 285358 337826 285410 337832
rect 285450 337884 285502 337890
rect 285450 337826 285502 337832
rect 285542 337884 285594 337890
rect 285632 337855 285688 337864
rect 285542 337826 285594 337832
rect 285048 337606 285122 337634
rect 285312 337680 285364 337686
rect 285312 337622 285364 337628
rect 285404 337680 285456 337686
rect 285456 337640 285536 337668
rect 285404 337622 285456 337628
rect 285048 337600 285076 337606
rect 284956 337572 285076 337600
rect 284852 334620 284904 334626
rect 284852 334562 284904 334568
rect 284852 326460 284904 326466
rect 284852 326402 284904 326408
rect 284760 326256 284812 326262
rect 284760 326198 284812 326204
rect 284760 326120 284812 326126
rect 284760 326062 284812 326068
rect 284668 171896 284720 171902
rect 284668 171838 284720 171844
rect 284772 171834 284800 326062
rect 284864 177682 284892 326402
rect 284852 177676 284904 177682
rect 284852 177618 284904 177624
rect 284956 177614 284984 337572
rect 285128 337544 285180 337550
rect 285128 337486 285180 337492
rect 285036 337476 285088 337482
rect 285036 337418 285088 337424
rect 285048 326126 285076 337418
rect 285140 326806 285168 337486
rect 285220 337476 285272 337482
rect 285220 337418 285272 337424
rect 285232 334801 285260 337418
rect 285324 336841 285352 337622
rect 285310 336832 285366 336841
rect 285310 336767 285366 336776
rect 285312 336592 285364 336598
rect 285312 336534 285364 336540
rect 285324 335481 285352 336534
rect 285508 335617 285536 337640
rect 285738 337600 285766 338028
rect 285830 337793 285858 338028
rect 285816 337784 285872 337793
rect 285816 337719 285872 337728
rect 285922 337668 285950 338028
rect 286014 337770 286042 338028
rect 286106 337890 286134 338028
rect 286198 337929 286226 338028
rect 286184 337920 286240 337929
rect 286094 337884 286146 337890
rect 286184 337855 286240 337864
rect 286094 337826 286146 337832
rect 286014 337742 286088 337770
rect 285922 337640 285996 337668
rect 285738 337572 285812 337600
rect 285588 337272 285640 337278
rect 285588 337214 285640 337220
rect 285600 336734 285628 337214
rect 285588 336728 285640 336734
rect 285588 336670 285640 336676
rect 285586 336424 285642 336433
rect 285586 336359 285642 336368
rect 285494 335608 285550 335617
rect 285494 335543 285550 335552
rect 285310 335472 285366 335481
rect 285310 335407 285366 335416
rect 285600 335034 285628 336359
rect 285784 336161 285812 337572
rect 285862 337512 285918 337521
rect 285862 337447 285918 337456
rect 285770 336152 285826 336161
rect 285770 336087 285826 336096
rect 285680 335368 285732 335374
rect 285680 335310 285732 335316
rect 285588 335028 285640 335034
rect 285588 334970 285640 334976
rect 285218 334792 285274 334801
rect 285218 334727 285274 334736
rect 285128 326800 285180 326806
rect 285128 326742 285180 326748
rect 285312 326732 285364 326738
rect 285312 326674 285364 326680
rect 285036 326120 285088 326126
rect 285036 326062 285088 326068
rect 284944 177608 284996 177614
rect 284944 177550 284996 177556
rect 284760 171828 284812 171834
rect 284760 171770 284812 171776
rect 284576 162240 284628 162246
rect 284576 162182 284628 162188
rect 284484 158092 284536 158098
rect 284484 158034 284536 158040
rect 284390 157992 284446 158001
rect 284390 157927 284446 157936
rect 285324 156670 285352 326674
rect 285692 326126 285720 335310
rect 285772 334076 285824 334082
rect 285772 334018 285824 334024
rect 285680 326120 285732 326126
rect 285680 326062 285732 326068
rect 285784 171134 285812 334018
rect 285876 173466 285904 337447
rect 285968 326262 285996 337640
rect 286060 326602 286088 337742
rect 286290 337736 286318 338028
rect 286382 337804 286410 338028
rect 286474 337958 286502 338028
rect 286566 337958 286594 338028
rect 286658 337958 286686 338028
rect 286462 337952 286514 337958
rect 286462 337894 286514 337900
rect 286554 337952 286606 337958
rect 286554 337894 286606 337900
rect 286646 337952 286698 337958
rect 286646 337894 286698 337900
rect 286508 337816 286560 337822
rect 286382 337776 286456 337804
rect 286290 337708 286364 337736
rect 286232 337612 286284 337618
rect 286232 337554 286284 337560
rect 286138 337512 286194 337521
rect 286138 337447 286194 337456
rect 286048 326596 286100 326602
rect 286048 326538 286100 326544
rect 286152 326346 286180 337447
rect 286244 334966 286272 337554
rect 286232 334960 286284 334966
rect 286232 334902 286284 334908
rect 286060 326318 286180 326346
rect 285956 326256 286008 326262
rect 285956 326198 286008 326204
rect 285956 326120 286008 326126
rect 285956 326062 286008 326068
rect 285864 173460 285916 173466
rect 285864 173402 285916 173408
rect 285968 173398 285996 326062
rect 286060 177478 286088 326318
rect 286140 326256 286192 326262
rect 286140 326198 286192 326204
rect 286152 177546 286180 326198
rect 286336 321554 286364 337708
rect 286428 335374 286456 337776
rect 286508 337758 286560 337764
rect 286600 337816 286652 337822
rect 286750 337793 286778 338028
rect 286842 337822 286870 338028
rect 286934 337963 286962 338028
rect 286920 337954 286976 337963
rect 287026 337958 287054 338028
rect 286920 337889 286976 337898
rect 287014 337952 287066 337958
rect 287014 337894 287066 337900
rect 286830 337816 286882 337822
rect 286600 337758 286652 337764
rect 286736 337784 286792 337793
rect 286416 335368 286468 335374
rect 286416 335310 286468 335316
rect 286520 332594 286548 337758
rect 286612 334082 286640 337758
rect 286830 337758 286882 337764
rect 286736 337719 286792 337728
rect 286692 337680 286744 337686
rect 286692 337622 286744 337628
rect 286876 337680 286928 337686
rect 287118 337668 287146 338028
rect 287210 337958 287238 338028
rect 287198 337952 287250 337958
rect 287302 337929 287330 338028
rect 287394 337958 287422 338028
rect 287486 337963 287514 338028
rect 287382 337952 287434 337958
rect 287198 337894 287250 337900
rect 287288 337920 287344 337929
rect 287382 337894 287434 337900
rect 287472 337954 287528 337963
rect 287578 337958 287606 338028
rect 287670 337958 287698 338028
rect 287762 337963 287790 338028
rect 287472 337889 287528 337898
rect 287566 337952 287618 337958
rect 287566 337894 287618 337900
rect 287658 337952 287710 337958
rect 287658 337894 287710 337900
rect 287748 337954 287804 337963
rect 287748 337889 287804 337898
rect 287288 337855 287344 337864
rect 287854 337822 287882 338028
rect 287946 337958 287974 338028
rect 288038 337958 288066 338028
rect 288130 337963 288158 338028
rect 287934 337952 287986 337958
rect 287934 337894 287986 337900
rect 288026 337952 288078 337958
rect 288026 337894 288078 337900
rect 288116 337954 288172 337963
rect 288222 337958 288250 338028
rect 288116 337889 288172 337898
rect 288210 337952 288262 337958
rect 288210 337894 288262 337900
rect 288314 337890 288342 338028
rect 288406 337963 288434 338028
rect 288392 337954 288448 337963
rect 288302 337884 288354 337890
rect 288392 337889 288448 337898
rect 288302 337826 288354 337832
rect 287244 337816 287296 337822
rect 287520 337816 287572 337822
rect 287244 337758 287296 337764
rect 287334 337784 287390 337793
rect 286876 337622 286928 337628
rect 287072 337640 287146 337668
rect 286704 334898 286732 337622
rect 286888 335209 286916 337622
rect 286968 337476 287020 337482
rect 286968 337418 287020 337424
rect 286874 335200 286930 335209
rect 286874 335135 286930 335144
rect 286692 334892 286744 334898
rect 286692 334834 286744 334840
rect 286600 334076 286652 334082
rect 286600 334018 286652 334024
rect 286428 332566 286548 332594
rect 286980 332594 287008 337418
rect 287072 336054 287100 337640
rect 287152 337544 287204 337550
rect 287152 337486 287204 337492
rect 287060 336048 287112 336054
rect 287060 335990 287112 335996
rect 286980 332566 287100 332594
rect 286428 326534 286456 332566
rect 286416 326528 286468 326534
rect 286416 326470 286468 326476
rect 286336 321526 286732 321554
rect 286140 177540 286192 177546
rect 286140 177482 286192 177488
rect 286048 177472 286100 177478
rect 286048 177414 286100 177420
rect 285956 173392 286008 173398
rect 285956 173334 286008 173340
rect 285784 171106 285904 171134
rect 285772 162172 285824 162178
rect 285772 162114 285824 162120
rect 285312 156664 285364 156670
rect 285312 156606 285364 156612
rect 285784 155924 285812 162114
rect 285876 159390 285904 171106
rect 286704 159458 286732 321526
rect 287072 160818 287100 332566
rect 287164 160886 287192 337486
rect 287256 336734 287284 337758
rect 287520 337758 287572 337764
rect 287842 337816 287894 337822
rect 288210 337816 288262 337822
rect 287842 337758 287894 337764
rect 288208 337784 288210 337793
rect 288262 337784 288264 337793
rect 287334 337719 287390 337728
rect 287244 336728 287296 336734
rect 287244 336670 287296 336676
rect 287244 336592 287296 336598
rect 287244 336534 287296 336540
rect 287256 335918 287284 336534
rect 287244 335912 287296 335918
rect 287244 335854 287296 335860
rect 287244 326392 287296 326398
rect 287244 326334 287296 326340
rect 287256 173330 287284 326334
rect 287348 174554 287376 337719
rect 287426 337648 287482 337657
rect 287426 337583 287482 337592
rect 287440 326398 287468 337583
rect 287428 326392 287480 326398
rect 287428 326334 287480 326340
rect 287428 326256 287480 326262
rect 287428 326198 287480 326204
rect 287440 177342 287468 326198
rect 287532 177410 287560 337758
rect 288498 337736 288526 338028
rect 288590 337958 288618 338028
rect 288578 337952 288630 337958
rect 288578 337894 288630 337900
rect 288682 337890 288710 338028
rect 288670 337884 288722 337890
rect 288670 337826 288722 337832
rect 288208 337719 288264 337728
rect 288360 337708 288526 337736
rect 288624 337748 288676 337754
rect 287612 337680 287664 337686
rect 287612 337622 287664 337628
rect 287796 337680 287848 337686
rect 287796 337622 287848 337628
rect 288256 337680 288308 337686
rect 288256 337622 288308 337628
rect 287624 337550 287652 337622
rect 287704 337612 287756 337618
rect 287704 337554 287756 337560
rect 287612 337544 287664 337550
rect 287612 337486 287664 337492
rect 287612 337408 287664 337414
rect 287612 337350 287664 337356
rect 287624 336666 287652 337350
rect 287612 336660 287664 336666
rect 287612 336602 287664 336608
rect 287610 336424 287666 336433
rect 287610 336359 287666 336368
rect 287624 336025 287652 336359
rect 287610 336016 287666 336025
rect 287610 335951 287666 335960
rect 287716 331214 287744 337554
rect 287624 331186 287744 331214
rect 287624 329118 287652 331186
rect 287612 329112 287664 329118
rect 287612 329054 287664 329060
rect 287808 326262 287836 337622
rect 288072 337612 288124 337618
rect 288072 337554 288124 337560
rect 288084 337464 288112 337554
rect 287992 337436 288112 337464
rect 287888 336524 287940 336530
rect 287888 336466 287940 336472
rect 287900 335918 287928 336466
rect 287888 335912 287940 335918
rect 287888 335854 287940 335860
rect 287796 326256 287848 326262
rect 287796 326198 287848 326204
rect 287992 316034 288020 337436
rect 288072 337340 288124 337346
rect 288072 337282 288124 337288
rect 288084 335714 288112 337282
rect 288072 335708 288124 335714
rect 288072 335650 288124 335656
rect 288268 334665 288296 337622
rect 288360 335374 288388 337708
rect 288624 337690 288676 337696
rect 288530 337512 288586 337521
rect 288440 337476 288492 337482
rect 288530 337447 288586 337456
rect 288440 337418 288492 337424
rect 288348 335368 288400 335374
rect 288348 335310 288400 335316
rect 288254 334656 288310 334665
rect 288254 334591 288310 334600
rect 287624 316006 288020 316034
rect 287624 193866 287652 316006
rect 287702 194576 287758 194585
rect 287702 194511 287758 194520
rect 287612 193860 287664 193866
rect 287612 193802 287664 193808
rect 287520 177404 287572 177410
rect 287520 177346 287572 177352
rect 287428 177336 287480 177342
rect 287428 177278 287480 177284
rect 287336 174548 287388 174554
rect 287336 174490 287388 174496
rect 287244 173324 287296 173330
rect 287244 173266 287296 173272
rect 287152 160880 287204 160886
rect 287152 160822 287204 160828
rect 287060 160812 287112 160818
rect 287060 160754 287112 160760
rect 286692 159452 286744 159458
rect 286692 159394 286744 159400
rect 285864 159384 285916 159390
rect 285864 159326 285916 159332
rect 287716 158030 287744 194511
rect 288452 160750 288480 337418
rect 288544 334540 288572 337447
rect 288636 334694 288664 337690
rect 288774 337634 288802 338028
rect 288866 337822 288894 338028
rect 288958 337963 288986 338028
rect 288944 337954 289000 337963
rect 288944 337889 289000 337898
rect 288854 337816 288906 337822
rect 289050 337770 289078 338028
rect 289142 337793 289170 338028
rect 289234 337958 289262 338028
rect 289222 337952 289274 337958
rect 289222 337894 289274 337900
rect 289326 337822 289354 338028
rect 289418 337822 289446 338028
rect 289314 337816 289366 337822
rect 288854 337758 288906 337764
rect 288958 337754 289078 337770
rect 288946 337748 289078 337754
rect 288998 337742 289078 337748
rect 289128 337784 289184 337793
rect 289314 337758 289366 337764
rect 289406 337816 289458 337822
rect 289510 337804 289538 338028
rect 289602 337963 289630 338028
rect 289588 337954 289644 337963
rect 289694 337958 289722 338028
rect 289786 337963 289814 338028
rect 289588 337889 289644 337898
rect 289682 337952 289734 337958
rect 289682 337894 289734 337900
rect 289772 337954 289828 337963
rect 289772 337889 289828 337898
rect 289878 337890 289906 338028
rect 289970 337890 289998 338028
rect 290062 337958 290090 338028
rect 290154 337963 290182 338028
rect 290050 337952 290102 337958
rect 290050 337894 290102 337900
rect 290140 337954 290196 337963
rect 290246 337958 290274 338028
rect 290338 337958 290366 338028
rect 290430 337963 290458 338028
rect 289866 337884 289918 337890
rect 289866 337826 289918 337832
rect 289958 337884 290010 337890
rect 290140 337889 290196 337898
rect 290234 337952 290286 337958
rect 290234 337894 290286 337900
rect 290326 337952 290378 337958
rect 290326 337894 290378 337900
rect 290416 337954 290472 337963
rect 290522 337958 290550 338028
rect 290628 338014 290780 338042
rect 290924 338030 290976 338036
rect 290416 337889 290472 337898
rect 290510 337952 290562 337958
rect 290510 337894 290562 337900
rect 289958 337826 290010 337832
rect 289510 337776 289584 337804
rect 289406 337758 289458 337764
rect 289128 337719 289184 337728
rect 288946 337690 288998 337696
rect 289176 337680 289228 337686
rect 288728 337606 288802 337634
rect 288898 337648 288954 337657
rect 288728 337249 288756 337606
rect 289176 337622 289228 337628
rect 288898 337583 288954 337592
rect 289084 337612 289136 337618
rect 288808 337544 288860 337550
rect 288808 337486 288860 337492
rect 288714 337240 288770 337249
rect 288714 337175 288770 337184
rect 288624 334688 288676 334694
rect 288624 334630 288676 334636
rect 288544 334512 288756 334540
rect 288532 334416 288584 334422
rect 288532 334358 288584 334364
rect 288544 162178 288572 334358
rect 288728 326777 288756 334512
rect 288714 326768 288770 326777
rect 288714 326703 288770 326712
rect 288820 326670 288848 337486
rect 288624 326664 288676 326670
rect 288624 326606 288676 326612
rect 288808 326664 288860 326670
rect 288808 326606 288860 326612
rect 288636 163538 288664 326606
rect 288714 326496 288770 326505
rect 288714 326431 288770 326440
rect 288728 173262 288756 326431
rect 288808 326392 288860 326398
rect 288808 326334 288860 326340
rect 288820 178838 288848 326334
rect 288912 178906 288940 337583
rect 289084 337554 289136 337560
rect 289096 331974 289124 337554
rect 289084 331968 289136 331974
rect 289084 331910 289136 331916
rect 289188 331906 289216 337622
rect 289360 337612 289412 337618
rect 289556 337600 289584 337776
rect 290278 337784 290334 337793
rect 289636 337748 289688 337754
rect 290096 337748 290148 337754
rect 289636 337690 289688 337696
rect 290016 337708 290096 337736
rect 289360 337554 289412 337560
rect 289464 337572 289584 337600
rect 289372 334422 289400 337554
rect 289360 334416 289412 334422
rect 289360 334358 289412 334364
rect 289176 331900 289228 331906
rect 289176 331842 289228 331848
rect 289464 326398 289492 337572
rect 289648 334626 289676 337690
rect 289728 337680 289780 337686
rect 289728 337622 289780 337628
rect 289912 337680 289964 337686
rect 289912 337622 289964 337628
rect 289740 335073 289768 337622
rect 289820 337612 289872 337618
rect 289820 337554 289872 337560
rect 289726 335064 289782 335073
rect 289726 334999 289782 335008
rect 289636 334620 289688 334626
rect 289636 334562 289688 334568
rect 289452 326392 289504 326398
rect 289452 326334 289504 326340
rect 289832 326346 289860 337554
rect 289924 326466 289952 337622
rect 289912 326460 289964 326466
rect 289912 326402 289964 326408
rect 289832 326318 289952 326346
rect 289820 326256 289872 326262
rect 289820 326198 289872 326204
rect 288900 178900 288952 178906
rect 288900 178842 288952 178848
rect 288808 178832 288860 178838
rect 288808 178774 288860 178780
rect 288716 173256 288768 173262
rect 288716 173198 288768 173204
rect 289832 167686 289860 326198
rect 289924 173194 289952 326318
rect 290016 178770 290044 337708
rect 290096 337690 290148 337696
rect 290200 337742 290278 337770
rect 290094 336696 290150 336705
rect 290094 336631 290150 336640
rect 290108 336161 290136 336631
rect 290094 336152 290150 336161
rect 290094 336087 290150 336096
rect 290200 327758 290228 337742
rect 290278 337719 290334 337728
rect 290372 337680 290424 337686
rect 290372 337622 290424 337628
rect 290464 337680 290516 337686
rect 290464 337622 290516 337628
rect 290384 332594 290412 337622
rect 290292 332566 290412 332594
rect 290188 327752 290240 327758
rect 290188 327694 290240 327700
rect 290292 321554 290320 332566
rect 290108 321526 290320 321554
rect 290004 178764 290056 178770
rect 290004 178706 290056 178712
rect 290108 178702 290136 321526
rect 290476 316034 290504 337622
rect 290646 335472 290702 335481
rect 290646 335407 290702 335416
rect 290660 321554 290688 335407
rect 290752 326262 290780 338014
rect 290832 338020 290884 338026
rect 290832 337962 290884 337968
rect 290844 330546 290872 337962
rect 290936 334830 290964 338030
rect 290924 334824 290976 334830
rect 290924 334766 290976 334772
rect 291028 334762 291056 338127
rect 293958 338056 294014 338065
rect 293958 337991 294014 338000
rect 292670 337920 292726 337929
rect 292670 337855 292726 337864
rect 291200 336728 291252 336734
rect 292684 336705 292712 337855
rect 292854 337240 292910 337249
rect 292854 337175 292910 337184
rect 292868 336802 292896 337175
rect 292856 336796 292908 336802
rect 292856 336738 292908 336744
rect 291200 336670 291252 336676
rect 292670 336696 292726 336705
rect 291016 334756 291068 334762
rect 291016 334698 291068 334704
rect 291212 332081 291240 336670
rect 292670 336631 292726 336640
rect 293408 336592 293460 336598
rect 293408 336534 293460 336540
rect 293224 336456 293276 336462
rect 293224 336398 293276 336404
rect 291936 336388 291988 336394
rect 291936 336330 291988 336336
rect 291844 335368 291896 335374
rect 291844 335310 291896 335316
rect 291198 332072 291254 332081
rect 291198 332007 291254 332016
rect 290832 330540 290884 330546
rect 290832 330482 290884 330488
rect 290740 326256 290792 326262
rect 290740 326198 290792 326204
rect 290660 321526 290780 321554
rect 290200 316006 290504 316034
rect 290200 180130 290228 316006
rect 290752 260166 290780 321526
rect 290740 260160 290792 260166
rect 290740 260102 290792 260108
rect 290188 180124 290240 180130
rect 290188 180066 290240 180072
rect 290096 178696 290148 178702
rect 290096 178638 290148 178644
rect 289912 173188 289964 173194
rect 289912 173130 289964 173136
rect 289820 167680 289872 167686
rect 289820 167622 289872 167628
rect 291856 166326 291884 335310
rect 291948 172378 291976 336330
rect 292120 335980 292172 335986
rect 292120 335922 292172 335928
rect 292028 335640 292080 335646
rect 292028 335582 292080 335588
rect 291936 172372 291988 172378
rect 291936 172314 291988 172320
rect 292040 172310 292068 335582
rect 292132 173534 292160 335922
rect 292120 173528 292172 173534
rect 292120 173470 292172 173476
rect 292028 172304 292080 172310
rect 292028 172246 292080 172252
rect 291844 166320 291896 166326
rect 291844 166262 291896 166268
rect 288624 163532 288676 163538
rect 288624 163474 288676 163480
rect 288532 162172 288584 162178
rect 288532 162114 288584 162120
rect 288440 160744 288492 160750
rect 288440 160686 288492 160692
rect 289634 158400 289690 158409
rect 289634 158335 289690 158344
rect 287704 158024 287756 158030
rect 287704 157966 287756 157972
rect 289648 155924 289676 158335
rect 293236 158098 293264 336398
rect 293316 335912 293368 335918
rect 293316 335854 293368 335860
rect 293328 166598 293356 335854
rect 293420 170746 293448 336534
rect 293500 335844 293552 335850
rect 293500 335786 293552 335792
rect 293512 176118 293540 335786
rect 293500 176112 293552 176118
rect 293500 176054 293552 176060
rect 293408 170740 293460 170746
rect 293408 170682 293460 170688
rect 293316 166592 293368 166598
rect 293316 166534 293368 166540
rect 293224 158092 293276 158098
rect 293224 158034 293276 158040
rect 293972 157418 294000 337991
rect 294604 335776 294656 335782
rect 294604 335718 294656 335724
rect 294512 326800 294564 326806
rect 294512 326742 294564 326748
rect 294524 326602 294552 326742
rect 294512 326596 294564 326602
rect 294512 326538 294564 326544
rect 294616 184278 294644 335718
rect 295982 335472 296038 335481
rect 295982 335407 296038 335416
rect 294604 184272 294656 184278
rect 294604 184214 294656 184220
rect 295996 172242 296024 335407
rect 296626 335336 296682 335345
rect 296626 335271 296682 335280
rect 296640 325825 296668 335271
rect 296626 325816 296682 325825
rect 296626 325751 296682 325760
rect 296626 325680 296682 325689
rect 296626 325615 296682 325624
rect 296640 316169 296668 325615
rect 296626 316160 296682 316169
rect 296626 316095 296682 316104
rect 296626 316024 296682 316033
rect 296626 315959 296682 315968
rect 296640 306513 296668 315959
rect 296626 306504 296682 306513
rect 296626 306439 296682 306448
rect 296626 306368 296682 306377
rect 296626 306303 296682 306312
rect 296640 296857 296668 306303
rect 296626 296848 296682 296857
rect 296626 296783 296682 296792
rect 296626 296712 296682 296721
rect 296626 296647 296682 296656
rect 296640 287201 296668 296647
rect 296626 287192 296682 287201
rect 296626 287127 296682 287136
rect 296626 287056 296682 287065
rect 296626 286991 296682 287000
rect 296640 277545 296668 286991
rect 296626 277536 296682 277545
rect 296626 277471 296682 277480
rect 296626 277400 296682 277409
rect 296626 277335 296682 277344
rect 296640 267889 296668 277335
rect 296626 267880 296682 267889
rect 296626 267815 296682 267824
rect 296626 267744 296682 267753
rect 296626 267679 296682 267688
rect 296640 248441 296668 267679
rect 296626 248432 296682 248441
rect 296626 248367 296682 248376
rect 296626 248296 296682 248305
rect 296626 248231 296682 248240
rect 296640 238785 296668 248231
rect 296626 238776 296682 238785
rect 296626 238711 296682 238720
rect 296626 238640 296682 238649
rect 296626 238575 296682 238584
rect 296640 229129 296668 238575
rect 296626 229120 296682 229129
rect 296626 229055 296682 229064
rect 296626 228984 296682 228993
rect 296626 228919 296682 228928
rect 296640 219473 296668 228919
rect 296626 219464 296682 219473
rect 296626 219399 296682 219408
rect 296626 219328 296682 219337
rect 296626 219263 296682 219272
rect 296640 209817 296668 219263
rect 296626 209808 296682 209817
rect 296626 209743 296682 209752
rect 296626 209672 296682 209681
rect 296626 209607 296682 209616
rect 296640 200161 296668 209607
rect 296626 200152 296682 200161
rect 296626 200087 296682 200096
rect 296626 200016 296682 200025
rect 296626 199951 296682 199960
rect 296640 190505 296668 199951
rect 296626 190496 296682 190505
rect 296626 190431 296682 190440
rect 296626 190360 296682 190369
rect 296626 190295 296682 190304
rect 296640 180849 296668 190295
rect 296626 180840 296682 180849
rect 296626 180775 296682 180784
rect 296626 180704 296682 180713
rect 296626 180639 296682 180648
rect 295984 172236 296036 172242
rect 295984 172178 296036 172184
rect 296640 171193 296668 180639
rect 296626 171184 296682 171193
rect 296626 171119 296682 171128
rect 296626 171048 296682 171057
rect 296626 170983 296682 170992
rect 296640 161537 296668 170983
rect 296626 161528 296682 161537
rect 296626 161463 296682 161472
rect 299492 161294 299520 382230
rect 299480 161288 299532 161294
rect 299480 161230 299532 161236
rect 298006 158672 298062 158681
rect 298006 158607 298062 158616
rect 293960 157412 294012 157418
rect 293960 157354 294012 157360
rect 293972 155938 294000 157354
rect 293972 155910 294170 155938
rect 298020 155924 298048 158607
rect 300136 157010 300164 384134
rect 300492 384124 300544 384130
rect 300492 384066 300544 384072
rect 300216 383852 300268 383858
rect 300216 383794 300268 383800
rect 300124 157004 300176 157010
rect 300124 156946 300176 156952
rect 300228 156942 300256 383794
rect 300400 383716 300452 383722
rect 300400 383658 300452 383664
rect 300308 382356 300360 382362
rect 300308 382298 300360 382304
rect 300320 157894 300348 382298
rect 300412 159594 300440 383658
rect 300504 262886 300532 384066
rect 301504 383784 301556 383790
rect 301504 383726 301556 383732
rect 300768 382696 300820 382702
rect 300768 382638 300820 382644
rect 300780 379506 300808 382638
rect 300952 381268 301004 381274
rect 300952 381210 301004 381216
rect 300860 381132 300912 381138
rect 300860 381074 300912 381080
rect 300768 379500 300820 379506
rect 300768 379442 300820 379448
rect 300492 262880 300544 262886
rect 300492 262822 300544 262828
rect 300400 159588 300452 159594
rect 300400 159530 300452 159536
rect 300872 158710 300900 381074
rect 300964 332246 300992 381210
rect 301042 380624 301098 380633
rect 301042 380559 301098 380568
rect 300952 332240 301004 332246
rect 300952 332182 301004 332188
rect 301056 332178 301084 380559
rect 301134 380488 301190 380497
rect 301134 380423 301190 380432
rect 301148 333606 301176 380423
rect 301136 333600 301188 333606
rect 301136 333542 301188 333548
rect 301044 332172 301096 332178
rect 301044 332114 301096 332120
rect 301516 158710 301544 383726
rect 301688 382832 301740 382838
rect 301688 382774 301740 382780
rect 301596 382424 301648 382430
rect 301596 382366 301648 382372
rect 300860 158704 300912 158710
rect 300860 158646 300912 158652
rect 301504 158704 301556 158710
rect 301504 158646 301556 158652
rect 300308 157888 300360 157894
rect 300308 157830 300360 157836
rect 301608 157826 301636 382366
rect 301700 157962 301728 382774
rect 301792 161401 301820 384270
rect 301884 302938 301912 384610
rect 343730 384432 343786 384441
rect 343730 384367 343786 384376
rect 322940 382968 322992 382974
rect 322940 382910 322992 382916
rect 306380 381676 306432 381682
rect 306380 381618 306432 381624
rect 301964 381200 302016 381206
rect 301964 381142 302016 381148
rect 301976 353258 302004 381142
rect 301964 353252 302016 353258
rect 301964 353194 302016 353200
rect 301872 302932 301924 302938
rect 301872 302874 301924 302880
rect 301778 161392 301834 161401
rect 301778 161327 301834 161336
rect 301688 157956 301740 157962
rect 301688 157898 301740 157904
rect 302514 157856 302570 157865
rect 301596 157820 301648 157826
rect 302514 157791 302570 157800
rect 301596 157762 301648 157768
rect 300216 156936 300268 156942
rect 300216 156878 300268 156884
rect 302528 155924 302556 157791
rect 306392 155924 306420 381618
rect 311162 336696 311218 336705
rect 311162 336631 311218 336640
rect 311176 163606 311204 336631
rect 311164 163600 311216 163606
rect 311164 163542 311216 163548
rect 310886 158536 310942 158545
rect 310886 158471 310942 158480
rect 310900 155924 310928 158471
rect 319260 157888 319312 157894
rect 319260 157830 319312 157836
rect 314752 157820 314804 157826
rect 314752 157762 314804 157768
rect 314764 155924 314792 157762
rect 319272 155924 319300 157830
rect 322952 155938 322980 382910
rect 337384 382628 337436 382634
rect 337384 382570 337436 382576
rect 335358 214568 335414 214577
rect 335358 214503 335414 214512
rect 335372 171134 335400 214503
rect 335372 171106 335584 171134
rect 327632 159588 327684 159594
rect 327632 159530 327684 159536
rect 322952 155910 323150 155938
rect 327644 155924 327672 159530
rect 331496 157956 331548 157962
rect 331496 157898 331548 157904
rect 331508 155924 331536 157898
rect 335556 155938 335584 171106
rect 337396 157962 337424 382570
rect 343638 158400 343694 158409
rect 343638 158335 343694 158344
rect 337384 157956 337436 157962
rect 337384 157898 337436 157904
rect 339868 157956 339920 157962
rect 339868 157898 339920 157904
rect 335556 155910 336030 155938
rect 339880 155924 339908 157898
rect 343652 155938 343680 158335
rect 343744 157457 343772 384367
rect 344652 384260 344704 384266
rect 344652 384202 344704 384208
rect 344284 384056 344336 384062
rect 344284 383998 344336 384004
rect 344100 383988 344152 383994
rect 344100 383930 344152 383936
rect 344008 381064 344060 381070
rect 344008 381006 344060 381012
rect 343916 337136 343968 337142
rect 343916 337078 343968 337084
rect 343730 157448 343786 157457
rect 343730 157383 343786 157392
rect 343652 155910 343758 155938
rect 284022 155680 284078 155689
rect 284022 155615 284078 155624
rect 271880 155382 271932 155388
rect 273166 155408 273222 155417
rect 269394 155343 269450 155352
rect 273166 155343 273222 155352
rect 259920 155236 259972 155242
rect 259920 155178 259972 155184
rect 342810 100736 342866 100745
rect 342866 100694 343114 100722
rect 342810 100671 342866 100680
rect 263692 100496 263744 100502
rect 263692 100438 263744 100444
rect 260840 100088 260892 100094
rect 260840 100030 260892 100036
rect 260024 97617 260052 100028
rect 260010 97608 260066 97617
rect 260010 97543 260066 97552
rect 260852 16574 260880 100030
rect 262220 100020 262272 100026
rect 262220 99962 262272 99968
rect 262232 16574 262260 99962
rect 263704 16574 263732 100438
rect 263888 97510 263916 100028
rect 267752 97986 267780 100028
rect 267740 97980 267792 97986
rect 267740 97922 267792 97928
rect 272260 97753 272288 100028
rect 276124 97782 276152 100028
rect 276112 97776 276164 97782
rect 272246 97744 272302 97753
rect 276112 97718 276164 97724
rect 272246 97679 272302 97688
rect 280632 97646 280660 100028
rect 284496 97714 284524 100028
rect 289004 97889 289032 100028
rect 288990 97880 289046 97889
rect 288990 97815 289046 97824
rect 284484 97708 284536 97714
rect 284484 97650 284536 97656
rect 280620 97640 280672 97646
rect 280620 97582 280672 97588
rect 292868 97578 292896 100028
rect 297376 97918 297404 100028
rect 297364 97912 297416 97918
rect 297364 97854 297416 97860
rect 301240 97850 301268 100028
rect 305012 100014 305762 100042
rect 301228 97844 301280 97850
rect 301228 97786 301280 97792
rect 292856 97572 292908 97578
rect 292856 97514 292908 97520
rect 263876 97504 263928 97510
rect 263876 97446 263928 97452
rect 305012 71738 305040 100014
rect 309612 97646 309640 100028
rect 309600 97640 309652 97646
rect 309600 97582 309652 97588
rect 314120 97578 314148 100028
rect 317984 97918 318012 100028
rect 317972 97912 318024 97918
rect 317972 97854 318024 97860
rect 322492 97782 322520 100028
rect 322480 97776 322532 97782
rect 322480 97718 322532 97724
rect 326356 97714 326384 100028
rect 330864 97889 330892 100028
rect 334728 97986 334756 100028
rect 334716 97980 334768 97986
rect 334716 97922 334768 97928
rect 330850 97880 330906 97889
rect 339236 97850 339264 100028
rect 330850 97815 330906 97824
rect 339224 97844 339276 97850
rect 339224 97786 339276 97792
rect 326344 97708 326396 97714
rect 326344 97650 326396 97656
rect 314108 97572 314160 97578
rect 314108 97514 314160 97520
rect 305000 71732 305052 71738
rect 305000 71674 305052 71680
rect 259840 16546 260696 16574
rect 260852 16546 261800 16574
rect 262232 16546 262536 16574
rect 263704 16546 264192 16574
rect 259472 6886 259684 6914
rect 259368 3664 259420 3670
rect 259368 3606 259420 3612
rect 259276 3256 259328 3262
rect 259276 3198 259328 3204
rect 259472 480 259500 6886
rect 260668 480 260696 16546
rect 261772 480 261800 16546
rect 258234 326 258488 354
rect 258234 -960 258346 326
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262508 354 262536 16546
rect 264164 480 264192 16546
rect 291384 9648 291436 9654
rect 291384 9590 291436 9596
rect 287796 9036 287848 9042
rect 287796 8978 287848 8984
rect 284300 8900 284352 8906
rect 284300 8842 284352 8848
rect 280712 8832 280764 8838
rect 280712 8774 280764 8780
rect 277124 8764 277176 8770
rect 277124 8706 277176 8712
rect 273628 6112 273680 6118
rect 273628 6054 273680 6060
rect 270040 6044 270092 6050
rect 270040 5986 270092 5992
rect 266544 5976 266596 5982
rect 266544 5918 266596 5924
rect 265348 3324 265400 3330
rect 265348 3266 265400 3272
rect 265360 480 265388 3266
rect 266556 480 266584 5918
rect 268844 4072 268896 4078
rect 268844 4014 268896 4020
rect 267740 3256 267792 3262
rect 267740 3198 267792 3204
rect 267752 480 267780 3198
rect 268856 480 268884 4014
rect 270052 480 270080 5986
rect 272432 4140 272484 4146
rect 272432 4082 272484 4088
rect 271236 3392 271288 3398
rect 271236 3334 271288 3340
rect 271248 480 271276 3334
rect 272444 480 272472 4082
rect 273640 480 273668 6054
rect 276020 3936 276072 3942
rect 274822 3904 274878 3913
rect 276020 3878 276072 3884
rect 274822 3839 274878 3848
rect 274836 480 274864 3839
rect 276032 480 276060 3878
rect 277136 480 277164 8706
rect 279516 6860 279568 6866
rect 279516 6802 279568 6808
rect 278320 3732 278372 3738
rect 278320 3674 278372 3680
rect 278332 480 278360 3674
rect 279528 480 279556 6802
rect 280724 480 280752 8774
rect 283104 6792 283156 6798
rect 283104 6734 283156 6740
rect 281908 4004 281960 4010
rect 281908 3946 281960 3952
rect 281920 480 281948 3946
rect 283116 480 283144 6734
rect 284312 480 284340 8842
rect 286600 6724 286652 6730
rect 286600 6666 286652 6672
rect 285404 3868 285456 3874
rect 285404 3810 285456 3816
rect 285416 480 285444 3810
rect 286612 480 286640 6666
rect 287808 480 287836 8978
rect 290188 6316 290240 6322
rect 290188 6258 290240 6264
rect 288992 3800 289044 3806
rect 288992 3742 289044 3748
rect 289004 480 289032 3742
rect 290200 480 290228 6258
rect 291396 480 291424 9590
rect 294880 9512 294932 9518
rect 294880 9454 294932 9460
rect 293684 6656 293736 6662
rect 293684 6598 293736 6604
rect 292580 3596 292632 3602
rect 292580 3538 292632 3544
rect 292592 480 292620 3538
rect 293696 480 293724 6598
rect 294892 480 294920 9454
rect 298468 9444 298520 9450
rect 298468 9386 298520 9392
rect 297272 6248 297324 6254
rect 297272 6190 297324 6196
rect 296076 3664 296128 3670
rect 296076 3606 296128 3612
rect 296088 480 296116 3606
rect 297284 480 297312 6190
rect 298480 480 298508 9386
rect 301964 9376 302016 9382
rect 301964 9318 302016 9324
rect 300768 6588 300820 6594
rect 300768 6530 300820 6536
rect 299664 3528 299716 3534
rect 299664 3470 299716 3476
rect 299676 480 299704 3470
rect 300780 480 300808 6530
rect 301976 480 302004 9318
rect 305552 9308 305604 9314
rect 305552 9250 305604 9256
rect 304356 6520 304408 6526
rect 304356 6462 304408 6468
rect 303160 3460 303212 3466
rect 303160 3402 303212 3408
rect 303172 480 303200 3402
rect 304368 480 304396 6462
rect 305564 480 305592 9250
rect 309048 9240 309100 9246
rect 309048 9182 309100 9188
rect 307944 6452 307996 6458
rect 307944 6394 307996 6400
rect 306746 3768 306802 3777
rect 306746 3703 306802 3712
rect 306760 480 306788 3703
rect 307956 480 307984 6394
rect 309060 480 309088 9182
rect 312636 9172 312688 9178
rect 312636 9114 312688 9120
rect 311440 6180 311492 6186
rect 311440 6122 311492 6128
rect 310242 3632 310298 3641
rect 310242 3567 310298 3576
rect 310256 480 310284 3567
rect 311452 480 311480 6122
rect 312648 480 312676 9114
rect 316224 8968 316276 8974
rect 316224 8910 316276 8916
rect 313830 3496 313886 3505
rect 313830 3431 313886 3440
rect 315028 3460 315080 3466
rect 313844 480 313872 3431
rect 315028 3402 315080 3408
rect 315040 480 315068 3402
rect 316236 480 316264 8910
rect 337476 6248 337528 6254
rect 337476 6190 337528 6196
rect 333888 6180 333940 6186
rect 333888 6122 333940 6128
rect 329196 4140 329248 4146
rect 329196 4082 329248 4088
rect 328000 4072 328052 4078
rect 328000 4014 328052 4020
rect 325608 4004 325660 4010
rect 325608 3946 325660 3952
rect 324412 3936 324464 3942
rect 324412 3878 324464 3884
rect 322112 3868 322164 3874
rect 322112 3810 322164 3816
rect 320916 3800 320968 3806
rect 320916 3742 320968 3748
rect 318524 3596 318576 3602
rect 318524 3538 318576 3544
rect 317326 3360 317382 3369
rect 317326 3295 317382 3304
rect 317340 480 317368 3295
rect 318536 480 318564 3538
rect 319720 3528 319772 3534
rect 319720 3470 319772 3476
rect 319732 480 319760 3470
rect 320928 480 320956 3742
rect 322124 480 322152 3810
rect 323308 3664 323360 3670
rect 323308 3606 323360 3612
rect 323320 480 323348 3606
rect 324424 480 324452 3878
rect 325620 480 325648 3946
rect 326804 3732 326856 3738
rect 326804 3674 326856 3680
rect 326816 480 326844 3674
rect 328012 480 328040 4014
rect 329208 480 329236 4082
rect 330392 3392 330444 3398
rect 330392 3334 330444 3340
rect 330404 480 330432 3334
rect 331588 3324 331640 3330
rect 331588 3266 331640 3272
rect 331600 480 331628 3266
rect 332692 3256 332744 3262
rect 332692 3198 332744 3204
rect 332704 480 332732 3198
rect 333900 480 333928 6122
rect 335082 3360 335138 3369
rect 335082 3295 335138 3304
rect 335096 480 335124 3295
rect 336278 3088 336334 3097
rect 336278 3023 336334 3032
rect 336292 480 336320 3023
rect 337488 480 337516 6190
rect 343362 3904 343418 3913
rect 343362 3839 343418 3848
rect 339866 3768 339922 3777
rect 339866 3703 339922 3712
rect 338670 3632 338726 3641
rect 338670 3567 338726 3576
rect 338684 480 338712 3567
rect 339880 480 339908 3703
rect 342166 3360 342222 3369
rect 342166 3295 342222 3304
rect 340970 3224 341026 3233
rect 340970 3159 341026 3168
rect 340984 480 341012 3159
rect 342180 480 342208 3295
rect 343376 480 343404 3839
rect 343928 3806 343956 337078
rect 344020 97578 344048 381006
rect 344112 103465 344140 383930
rect 344192 155576 344244 155582
rect 344192 155518 344244 155524
rect 344098 103456 344154 103465
rect 344098 103391 344154 103400
rect 344008 97572 344060 97578
rect 344008 97514 344060 97520
rect 344204 4049 344232 155518
rect 344296 130422 344324 383998
rect 344376 155508 344428 155514
rect 344376 155450 344428 155456
rect 344284 130416 344336 130422
rect 344284 130358 344336 130364
rect 344190 4040 344246 4049
rect 344388 4010 344416 155450
rect 344468 155440 344520 155446
rect 344468 155382 344520 155388
rect 344190 3975 344246 3984
rect 344376 4004 344428 4010
rect 344376 3946 344428 3952
rect 343916 3800 343968 3806
rect 343916 3742 343968 3748
rect 344480 3641 344508 155382
rect 344560 155372 344612 155378
rect 344560 155314 344612 155320
rect 344572 16574 344600 155314
rect 344664 151745 344692 384202
rect 523682 384160 523738 384169
rect 523682 384095 523738 384104
rect 347780 383920 347832 383926
rect 347780 383862 347832 383868
rect 347042 381712 347098 381721
rect 347042 381647 347098 381656
rect 346584 337408 346636 337414
rect 346584 337350 346636 337356
rect 345664 337272 345716 337278
rect 345664 337214 345716 337220
rect 345112 302932 345164 302938
rect 345112 302874 345164 302880
rect 345020 157004 345072 157010
rect 345020 156946 345072 156952
rect 344650 151736 344706 151745
rect 344650 151671 344706 151680
rect 344650 148336 344706 148345
rect 344650 148271 344706 148280
rect 344664 97646 344692 148271
rect 345032 134065 345060 156946
rect 345124 147665 345152 302874
rect 345204 262880 345256 262886
rect 345204 262822 345256 262828
rect 345110 147656 345166 147665
rect 345110 147591 345166 147600
rect 345018 134056 345074 134065
rect 345018 133991 345074 134000
rect 345020 130416 345072 130422
rect 345020 130358 345072 130364
rect 344926 129840 344982 129849
rect 344926 129775 344982 129784
rect 344652 97640 344704 97646
rect 344652 97582 344704 97588
rect 344572 16546 344692 16574
rect 344466 3632 344522 3641
rect 344664 3602 344692 16546
rect 344940 6866 344968 129775
rect 345032 116385 345060 130358
rect 345018 116376 345074 116385
rect 345018 116311 345074 116320
rect 345216 107545 345244 262822
rect 345386 180024 345442 180033
rect 345386 179959 345442 179968
rect 345294 158264 345350 158273
rect 345294 158199 345350 158208
rect 345202 107536 345258 107545
rect 345202 107471 345258 107480
rect 344928 6860 344980 6866
rect 344928 6802 344980 6808
rect 344834 3632 344890 3641
rect 344466 3567 344522 3576
rect 344652 3596 344704 3602
rect 344834 3567 344890 3576
rect 344652 3538 344704 3544
rect 344558 3496 344614 3505
rect 344558 3431 344614 3440
rect 344572 480 344600 3431
rect 344848 3233 344876 3567
rect 345308 3505 345336 158199
rect 345400 112305 345428 179959
rect 345478 170504 345534 170513
rect 345478 170439 345534 170448
rect 345492 125225 345520 170439
rect 345572 158704 345624 158710
rect 345572 158646 345624 158652
rect 345584 129985 345612 158646
rect 345570 129976 345626 129985
rect 345570 129911 345626 129920
rect 345478 125216 345534 125225
rect 345478 125151 345534 125160
rect 345386 112296 345442 112305
rect 345386 112231 345442 112240
rect 345676 16574 345704 337214
rect 346492 337204 346544 337210
rect 346492 337146 346544 337152
rect 346400 337068 346452 337074
rect 346400 337010 346452 337016
rect 345756 156936 345808 156942
rect 345756 156878 345808 156884
rect 345768 138825 345796 156878
rect 345846 155544 345902 155553
rect 345846 155479 345902 155488
rect 345754 138816 345810 138825
rect 345754 138751 345810 138760
rect 345676 16546 345796 16574
rect 345294 3496 345350 3505
rect 345294 3431 345350 3440
rect 344834 3224 344890 3233
rect 344834 3159 344890 3168
rect 345768 480 345796 16546
rect 345860 3874 345888 155479
rect 345848 3868 345900 3874
rect 345848 3810 345900 3816
rect 346412 3466 346440 337010
rect 346400 3460 346452 3466
rect 346400 3402 346452 3408
rect 346504 3369 346532 337146
rect 346490 3360 346546 3369
rect 346596 3330 346624 337350
rect 346676 337340 346728 337346
rect 346676 337282 346728 337288
rect 346688 4078 346716 337282
rect 346768 336320 346820 336326
rect 346768 336262 346820 336268
rect 346676 4072 346728 4078
rect 346676 4014 346728 4020
rect 346780 3942 346808 336262
rect 346860 335300 346912 335306
rect 346860 335242 346912 335248
rect 346768 3936 346820 3942
rect 346768 3878 346820 3884
rect 346490 3295 346546 3304
rect 346584 3324 346636 3330
rect 346584 3266 346636 3272
rect 346872 3262 346900 335242
rect 346952 158636 347004 158642
rect 346952 158578 347004 158584
rect 346860 3256 346912 3262
rect 346860 3198 346912 3204
rect 346964 480 346992 158578
rect 347056 126954 347084 381647
rect 347136 155304 347188 155310
rect 347136 155246 347188 155252
rect 347044 126948 347096 126954
rect 347044 126890 347096 126896
rect 347148 3097 347176 155246
rect 347228 155236 347280 155242
rect 347228 155178 347280 155184
rect 347240 4146 347268 155178
rect 347792 97782 347820 383862
rect 356702 383752 356758 383761
rect 356702 383687 356758 383696
rect 349252 382560 349304 382566
rect 349252 382502 349304 382508
rect 347872 382492 347924 382498
rect 347872 382434 347924 382440
rect 347884 97850 347912 382434
rect 349160 335232 349212 335238
rect 349160 335174 349212 335180
rect 348330 161256 348386 161265
rect 347964 161220 348016 161226
rect 348330 161191 348386 161200
rect 347964 161162 348016 161168
rect 347872 97844 347924 97850
rect 347872 97786 347924 97792
rect 347780 97776 347832 97782
rect 347780 97718 347832 97724
rect 347976 11898 348004 161162
rect 348240 161152 348292 161158
rect 348240 161094 348292 161100
rect 348056 158568 348108 158574
rect 348056 158510 348108 158516
rect 347964 11892 348016 11898
rect 347964 11834 348016 11840
rect 348068 11778 348096 158510
rect 348146 158128 348202 158137
rect 348146 158063 348202 158072
rect 347884 11750 348096 11778
rect 347228 4140 347280 4146
rect 347228 4082 347280 4088
rect 347884 3398 347912 11750
rect 348056 11688 348108 11694
rect 348056 11630 348108 11636
rect 347872 3392 347924 3398
rect 347872 3334 347924 3340
rect 347134 3088 347190 3097
rect 347134 3023 347190 3032
rect 348068 480 348096 11630
rect 348160 3670 348188 158063
rect 348252 6254 348280 161094
rect 348344 97714 348372 161191
rect 348332 97708 348384 97714
rect 348332 97650 348384 97656
rect 349172 16574 349200 335174
rect 349264 97918 349292 382502
rect 351920 335164 351972 335170
rect 351920 335106 351972 335112
rect 349344 169244 349396 169250
rect 349344 169186 349396 169192
rect 349252 97912 349304 97918
rect 349252 97854 349304 97860
rect 349172 16546 349292 16574
rect 348240 6248 348292 6254
rect 348240 6190 348292 6196
rect 348148 3664 348200 3670
rect 348148 3606 348200 3612
rect 349264 480 349292 16546
rect 349356 3482 349384 169186
rect 350540 161084 350592 161090
rect 350540 161026 350592 161032
rect 349434 160984 349490 160993
rect 349434 160919 349490 160928
rect 349448 3641 349476 160919
rect 349712 158500 349764 158506
rect 349712 158442 349764 158448
rect 349528 158432 349580 158438
rect 349528 158374 349580 158380
rect 349540 3738 349568 158374
rect 349620 158296 349672 158302
rect 349620 158238 349672 158244
rect 349528 3732 349580 3738
rect 349528 3674 349580 3680
rect 349434 3632 349490 3641
rect 349632 3602 349660 158238
rect 349724 3777 349752 158442
rect 349804 158364 349856 158370
rect 349804 158306 349856 158312
rect 349816 6186 349844 158306
rect 349894 155680 349950 155689
rect 349894 155615 349950 155624
rect 349908 97986 349936 155615
rect 349896 97980 349948 97986
rect 349896 97922 349948 97928
rect 350552 16574 350580 161026
rect 351932 16574 351960 335106
rect 354680 332104 354732 332110
rect 354680 332046 354732 332052
rect 353300 158228 353352 158234
rect 353300 158170 353352 158176
rect 353312 16574 353340 158170
rect 354692 16574 354720 332046
rect 356058 155408 356114 155417
rect 356058 155343 356114 155352
rect 356072 16574 356100 155343
rect 350552 16546 351224 16574
rect 351932 16546 352880 16574
rect 353312 16546 353616 16574
rect 354692 16546 355272 16574
rect 356072 16546 356376 16574
rect 349804 6180 349856 6186
rect 349804 6122 349856 6128
rect 349710 3768 349766 3777
rect 349710 3703 349766 3712
rect 349434 3567 349490 3576
rect 349620 3596 349672 3602
rect 349620 3538 349672 3544
rect 349356 3454 350488 3482
rect 350460 480 350488 3454
rect 262926 354 263038 480
rect 262508 326 263038 354
rect 262926 -960 263038 326
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351196 354 351224 16546
rect 352852 480 352880 16546
rect 351614 354 351726 480
rect 351196 326 351726 354
rect 351614 -960 351726 326
rect 352810 -960 352922 480
rect 353588 354 353616 16546
rect 355244 480 355272 16546
rect 356348 480 356376 16546
rect 356716 3466 356744 383687
rect 407762 381304 407818 381313
rect 407762 381239 407818 381248
rect 394700 337000 394752 337006
rect 394700 336942 394752 336948
rect 382922 336560 382978 336569
rect 382922 336495 382978 336504
rect 379520 332036 379572 332042
rect 379520 331978 379572 331984
rect 361580 330676 361632 330682
rect 361580 330618 361632 330624
rect 358820 330608 358872 330614
rect 358820 330550 358872 330556
rect 357440 163736 357492 163742
rect 357440 163678 357492 163684
rect 356704 3460 356756 3466
rect 356704 3402 356756 3408
rect 357452 2242 357480 163678
rect 357532 158160 357584 158166
rect 357532 158102 357584 158108
rect 357440 2236 357492 2242
rect 357440 2178 357492 2184
rect 357544 480 357572 158102
rect 358832 16574 358860 330550
rect 360200 156868 360252 156874
rect 360200 156810 360252 156816
rect 360212 16574 360240 156810
rect 361592 16574 361620 330618
rect 365720 326664 365772 326670
rect 365720 326606 365772 326612
rect 364340 170808 364392 170814
rect 364340 170750 364392 170756
rect 362960 163940 363012 163946
rect 362960 163882 363012 163888
rect 362972 16574 363000 163882
rect 364352 16574 364380 170750
rect 358832 16546 359504 16574
rect 360212 16546 361160 16574
rect 361592 16546 361896 16574
rect 362972 16546 363552 16574
rect 364352 16546 364656 16574
rect 358728 2236 358780 2242
rect 358728 2178 358780 2184
rect 358740 480 358768 2178
rect 354006 354 354118 480
rect 353588 326 354118 354
rect 354006 -960 354118 326
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359476 354 359504 16546
rect 361132 480 361160 16546
rect 359894 354 360006 480
rect 359476 326 360006 354
rect 359894 -960 360006 326
rect 361090 -960 361202 480
rect 361868 354 361896 16546
rect 363524 480 363552 16546
rect 364628 480 364656 16546
rect 365732 3346 365760 326606
rect 376760 325032 376812 325038
rect 376760 324974 376812 324980
rect 373998 320784 374054 320793
rect 373998 320719 374054 320728
rect 368480 179104 368532 179110
rect 368480 179046 368532 179052
rect 367100 174820 367152 174826
rect 367100 174762 367152 174768
rect 365812 163872 365864 163878
rect 365812 163814 365864 163820
rect 365824 3534 365852 163814
rect 367112 16574 367140 174762
rect 368492 16574 368520 179046
rect 371240 174752 371292 174758
rect 371240 174694 371292 174700
rect 369860 163804 369912 163810
rect 369860 163746 369912 163752
rect 369872 16574 369900 163746
rect 367112 16546 367784 16574
rect 368492 16546 369440 16574
rect 369872 16546 370176 16574
rect 365812 3528 365864 3534
rect 365812 3470 365864 3476
rect 367008 3528 367060 3534
rect 367008 3470 367060 3476
rect 365732 3318 365852 3346
rect 365824 480 365852 3318
rect 367020 480 367048 3470
rect 362286 354 362398 480
rect 361868 326 362398 354
rect 362286 -960 362398 326
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 367756 354 367784 16546
rect 369412 480 369440 16546
rect 368174 354 368286 480
rect 367756 326 368286 354
rect 368174 -960 368286 326
rect 369370 -960 369482 480
rect 370148 354 370176 16546
rect 370566 354 370678 480
rect 370148 326 370678 354
rect 371252 354 371280 174694
rect 372620 162308 372672 162314
rect 372620 162250 372672 162256
rect 372632 16574 372660 162250
rect 372632 16546 372936 16574
rect 372908 480 372936 16546
rect 374012 3346 374040 320719
rect 374090 174720 374146 174729
rect 374090 174655 374146 174664
rect 374104 3534 374132 174655
rect 375378 165064 375434 165073
rect 375378 164999 375434 165008
rect 375392 16574 375420 164999
rect 376772 16574 376800 324974
rect 378140 174684 378192 174690
rect 378140 174626 378192 174632
rect 378152 16574 378180 174626
rect 375392 16546 376064 16574
rect 376772 16546 377720 16574
rect 378152 16546 378456 16574
rect 374092 3528 374144 3534
rect 374092 3470 374144 3476
rect 375288 3528 375340 3534
rect 375288 3470 375340 3476
rect 374012 3318 374132 3346
rect 374104 480 374132 3318
rect 375300 480 375328 3470
rect 371670 354 371782 480
rect 371252 326 371782 354
rect 370566 -960 370678 326
rect 371670 -960 371782 326
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376036 354 376064 16546
rect 377692 480 377720 16546
rect 376454 354 376566 480
rect 376036 326 376566 354
rect 376454 -960 376566 326
rect 377650 -960 377762 480
rect 378428 354 378456 16546
rect 378846 354 378958 480
rect 378428 326 378958 354
rect 379532 354 379560 331978
rect 382280 176452 382332 176458
rect 382280 176394 382332 176400
rect 380900 163668 380952 163674
rect 380900 163610 380952 163616
rect 380912 16574 380940 163610
rect 380912 16546 381216 16574
rect 381188 480 381216 16546
rect 382292 3346 382320 176394
rect 382372 165300 382424 165306
rect 382372 165242 382424 165248
rect 382384 3534 382412 165242
rect 382936 159594 382964 336495
rect 391938 333704 391994 333713
rect 391938 333639 391994 333648
rect 386420 179036 386472 179042
rect 386420 178978 386472 178984
rect 385040 176384 385092 176390
rect 385040 176326 385092 176332
rect 383660 165232 383712 165238
rect 383660 165174 383712 165180
rect 382924 159588 382976 159594
rect 382924 159530 382976 159536
rect 383672 16574 383700 165174
rect 385052 16574 385080 176326
rect 386432 16574 386460 178978
rect 389180 176316 389232 176322
rect 389180 176258 389232 176264
rect 387800 165164 387852 165170
rect 387800 165106 387852 165112
rect 383672 16546 384344 16574
rect 385052 16546 386000 16574
rect 386432 16546 386736 16574
rect 382372 3528 382424 3534
rect 382372 3470 382424 3476
rect 383568 3528 383620 3534
rect 383568 3470 383620 3476
rect 382292 3318 382412 3346
rect 382384 480 382412 3318
rect 383580 480 383608 3470
rect 379950 354 380062 480
rect 379532 326 380062 354
rect 378846 -960 378958 326
rect 379950 -960 380062 326
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384316 354 384344 16546
rect 385972 480 386000 16546
rect 384734 354 384846 480
rect 384316 326 384846 354
rect 384734 -960 384846 326
rect 385930 -960 386042 480
rect 386708 354 386736 16546
rect 387126 354 387238 480
rect 386708 326 387238 354
rect 387812 354 387840 165106
rect 389192 16574 389220 176258
rect 390652 165096 390704 165102
rect 390652 165038 390704 165044
rect 390558 164928 390614 164937
rect 390558 164863 390614 164872
rect 389192 16546 389496 16574
rect 389468 480 389496 16546
rect 390572 3346 390600 164863
rect 390664 3534 390692 165038
rect 391952 16574 391980 333639
rect 393320 172372 393372 172378
rect 393320 172314 393372 172320
rect 393332 16574 393360 172314
rect 394712 16574 394740 336942
rect 398840 333532 398892 333538
rect 398840 333474 398892 333480
rect 396080 323604 396132 323610
rect 396080 323546 396132 323552
rect 391952 16546 392624 16574
rect 393332 16546 394280 16574
rect 394712 16546 395384 16574
rect 390652 3528 390704 3534
rect 390652 3470 390704 3476
rect 391848 3528 391900 3534
rect 391848 3470 391900 3476
rect 390572 3318 390692 3346
rect 390664 480 390692 3318
rect 391860 480 391888 3470
rect 388230 354 388342 480
rect 387812 326 388342 354
rect 387126 -960 387238 326
rect 388230 -960 388342 326
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 392596 354 392624 16546
rect 394252 480 394280 16546
rect 395356 480 395384 16546
rect 393014 354 393126 480
rect 392596 326 393126 354
rect 393014 -960 393126 326
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396092 354 396120 323546
rect 397460 172304 397512 172310
rect 397460 172246 397512 172252
rect 397472 16574 397500 172246
rect 397472 16546 397776 16574
rect 397748 480 397776 16546
rect 398852 2242 398880 333474
rect 407120 333464 407172 333470
rect 407120 333406 407172 333412
rect 398932 327888 398984 327894
rect 398932 327830 398984 327836
rect 398840 2236 398892 2242
rect 398840 2178 398892 2184
rect 398944 480 398972 327830
rect 402980 176248 403032 176254
rect 402980 176190 403032 176196
rect 400220 165028 400272 165034
rect 400220 164970 400272 164976
rect 400232 16574 400260 164970
rect 401600 164960 401652 164966
rect 401600 164902 401652 164908
rect 401612 16574 401640 164902
rect 402992 16574 403020 176190
rect 404360 173528 404412 173534
rect 404360 173470 404412 173476
rect 400232 16546 400904 16574
rect 401612 16546 402560 16574
rect 402992 16546 403664 16574
rect 400128 2236 400180 2242
rect 400128 2178 400180 2184
rect 400140 480 400168 2178
rect 396510 354 396622 480
rect 396092 326 396622 354
rect 396510 -960 396622 326
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 400876 354 400904 16546
rect 402532 480 402560 16546
rect 403636 480 403664 16546
rect 401294 354 401406 480
rect 400876 326 401406 354
rect 401294 -960 401406 326
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404372 354 404400 173470
rect 405740 164892 405792 164898
rect 405740 164834 405792 164840
rect 405752 16574 405780 164834
rect 405752 16546 406056 16574
rect 406028 480 406056 16546
rect 407132 3346 407160 333406
rect 407210 175944 407266 175953
rect 407210 175879 407266 175888
rect 407224 3534 407252 175879
rect 407776 167006 407804 381239
rect 430580 338292 430632 338298
rect 430580 338234 430632 338240
rect 408500 336932 408552 336938
rect 408500 336874 408552 336880
rect 407764 167000 407816 167006
rect 407764 166942 407816 166948
rect 408512 16574 408540 336874
rect 427818 333568 427874 333577
rect 427818 333503 427874 333512
rect 414020 333396 414072 333402
rect 414020 333338 414072 333344
rect 412640 166660 412692 166666
rect 412640 166602 412692 166608
rect 409878 159624 409934 159633
rect 409878 159559 409934 159568
rect 409892 16574 409920 159559
rect 411260 158092 411312 158098
rect 411260 158034 411312 158040
rect 411272 16574 411300 158034
rect 408512 16546 409184 16574
rect 409892 16546 410840 16574
rect 411272 16546 411944 16574
rect 407212 3528 407264 3534
rect 407212 3470 407264 3476
rect 408408 3528 408460 3534
rect 408408 3470 408460 3476
rect 407132 3318 407252 3346
rect 407224 480 407252 3318
rect 408420 480 408448 3470
rect 404790 354 404902 480
rect 404372 326 404902 354
rect 404790 -960 404902 326
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409156 354 409184 16546
rect 410812 480 410840 16546
rect 411916 480 411944 16546
rect 409574 354 409686 480
rect 409156 326 409686 354
rect 409574 -960 409686 326
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 412652 354 412680 166602
rect 414032 16574 414060 333338
rect 420920 333328 420972 333334
rect 420920 333270 420972 333276
rect 418160 180192 418212 180198
rect 418160 180134 418212 180140
rect 415400 178968 415452 178974
rect 415400 178910 415452 178916
rect 414032 16546 414336 16574
rect 414308 480 414336 16546
rect 415412 3346 415440 178910
rect 416780 176180 416832 176186
rect 416780 176122 416832 176128
rect 415492 166524 415544 166530
rect 415492 166466 415544 166472
rect 415504 3534 415532 166466
rect 416792 16574 416820 176122
rect 418172 16574 418200 180134
rect 419540 166456 419592 166462
rect 419540 166398 419592 166404
rect 419552 16574 419580 166398
rect 416792 16546 417464 16574
rect 418172 16546 418568 16574
rect 419552 16546 420224 16574
rect 415492 3528 415544 3534
rect 415492 3470 415544 3476
rect 416688 3528 416740 3534
rect 416688 3470 416740 3476
rect 415412 3318 415532 3346
rect 415504 480 415532 3318
rect 416700 480 416728 3470
rect 413070 354 413182 480
rect 412652 326 413182 354
rect 413070 -960 413182 326
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417436 354 417464 16546
rect 417854 354 417966 480
rect 417436 326 417966 354
rect 418540 354 418568 16546
rect 420196 480 420224 16546
rect 418958 354 419070 480
rect 418540 326 419070 354
rect 417854 -960 417966 326
rect 418958 -960 419070 326
rect 420154 -960 420266 480
rect 420932 354 420960 333270
rect 423680 327820 423732 327826
rect 423680 327762 423732 327768
rect 422300 170740 422352 170746
rect 422300 170682 422352 170688
rect 422312 16574 422340 170682
rect 422312 16546 422616 16574
rect 422588 480 422616 16546
rect 423692 3346 423720 327762
rect 423772 176044 423824 176050
rect 423772 175986 423824 175992
rect 423784 3534 423812 175986
rect 425058 166560 425114 166569
rect 425058 166495 425114 166504
rect 425072 16574 425100 166495
rect 426438 166424 426494 166433
rect 426438 166359 426494 166368
rect 426452 16574 426480 166359
rect 427832 16574 427860 333503
rect 429200 166592 429252 166598
rect 429200 166534 429252 166540
rect 425072 16546 425744 16574
rect 426452 16546 426848 16574
rect 427832 16546 428504 16574
rect 423772 3528 423824 3534
rect 423772 3470 423824 3476
rect 424968 3528 425020 3534
rect 424968 3470 425020 3476
rect 423692 3318 423812 3346
rect 423784 480 423812 3318
rect 424980 480 425008 3470
rect 421350 354 421462 480
rect 420932 326 421462 354
rect 421350 -960 421462 326
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 425716 354 425744 16546
rect 426134 354 426246 480
rect 425716 326 426246 354
rect 426820 354 426848 16546
rect 428476 480 428504 16546
rect 427238 354 427350 480
rect 426820 326 427350 354
rect 426134 -960 426246 326
rect 427238 -960 427350 326
rect 428434 -960 428546 480
rect 429212 354 429240 166534
rect 430592 16574 430620 338234
rect 448520 338224 448572 338230
rect 448520 338166 448572 338172
rect 445758 333432 445814 333441
rect 445758 333367 445814 333376
rect 438860 333260 438912 333266
rect 438860 333202 438912 333208
rect 436100 176112 436152 176118
rect 436100 176054 436152 176060
rect 431960 175976 432012 175982
rect 431960 175918 432012 175924
rect 430592 16546 430896 16574
rect 430868 480 430896 16546
rect 431972 3346 432000 175918
rect 432052 170672 432104 170678
rect 432052 170614 432104 170620
rect 432064 3534 432092 170614
rect 434720 170604 434772 170610
rect 434720 170546 434772 170552
rect 433340 168156 433392 168162
rect 433340 168098 433392 168104
rect 433352 16574 433380 168098
rect 434732 16574 434760 170546
rect 436112 16574 436140 176054
rect 437480 168088 437532 168094
rect 437480 168030 437532 168036
rect 433352 16546 434024 16574
rect 434732 16546 435128 16574
rect 436112 16546 436784 16574
rect 432052 3528 432104 3534
rect 432052 3470 432104 3476
rect 433248 3528 433300 3534
rect 433248 3470 433300 3476
rect 431972 3318 432092 3346
rect 432064 480 432092 3318
rect 433260 480 433288 3470
rect 429630 354 429742 480
rect 429212 326 429742 354
rect 429630 -960 429742 326
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 433996 354 434024 16546
rect 434414 354 434526 480
rect 433996 326 434526 354
rect 435100 354 435128 16546
rect 436756 480 436784 16546
rect 435518 354 435630 480
rect 435100 326 435630 354
rect 434414 -960 434526 326
rect 435518 -960 435630 326
rect 436714 -960 436826 480
rect 437492 354 437520 168030
rect 438872 16574 438900 333202
rect 443000 260160 443052 260166
rect 443000 260102 443052 260108
rect 441620 170536 441672 170542
rect 441620 170478 441672 170484
rect 440240 168020 440292 168026
rect 440240 167962 440292 167968
rect 438872 16546 439176 16574
rect 439148 480 439176 16546
rect 440252 2242 440280 167962
rect 440332 166388 440384 166394
rect 440332 166330 440384 166336
rect 440240 2236 440292 2242
rect 440240 2178 440292 2184
rect 440344 480 440372 166330
rect 441632 16574 441660 170478
rect 443012 16574 443040 260102
rect 444378 186960 444434 186969
rect 444378 186895 444434 186904
rect 444392 16574 444420 186895
rect 441632 16546 442672 16574
rect 443012 16546 443408 16574
rect 444392 16546 445064 16574
rect 441528 2236 441580 2242
rect 441528 2178 441580 2184
rect 441540 480 441568 2178
rect 442644 480 442672 16546
rect 437910 354 438022 480
rect 437492 326 438022 354
rect 437910 -960 438022 326
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443380 354 443408 16546
rect 445036 480 445064 16546
rect 443798 354 443910 480
rect 443380 326 443910 354
rect 443798 -960 443910 326
rect 444994 -960 445106 480
rect 445772 354 445800 333367
rect 447138 166288 447194 166297
rect 447138 166223 447194 166232
rect 447152 16574 447180 166223
rect 447152 16546 447456 16574
rect 447428 480 447456 16546
rect 448532 3346 448560 338166
rect 465080 338156 465132 338162
rect 465080 338098 465132 338104
rect 451280 336864 451332 336870
rect 451280 336806 451332 336812
rect 449900 184272 449952 184278
rect 449900 184214 449952 184220
rect 448612 161016 448664 161022
rect 448612 160958 448664 160964
rect 448624 3534 448652 160958
rect 449912 16574 449940 184214
rect 451292 16574 451320 336806
rect 463698 333296 463754 333305
rect 463698 333231 463754 333240
rect 456800 324964 456852 324970
rect 456800 324906 456852 324912
rect 452660 177812 452712 177818
rect 452660 177754 452712 177760
rect 452672 16574 452700 177754
rect 454040 174616 454092 174622
rect 454040 174558 454092 174564
rect 449912 16546 450952 16574
rect 451292 16546 451688 16574
rect 452672 16546 453344 16574
rect 448612 3528 448664 3534
rect 448612 3470 448664 3476
rect 449808 3528 449860 3534
rect 449808 3470 449860 3476
rect 448532 3318 448652 3346
rect 448624 480 448652 3318
rect 449820 480 449848 3470
rect 450924 480 450952 16546
rect 446190 354 446302 480
rect 445772 326 446302 354
rect 446190 -960 446302 326
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 451660 354 451688 16546
rect 453316 480 453344 16546
rect 452078 354 452190 480
rect 451660 326 452190 354
rect 452078 -960 452190 326
rect 453274 -960 453386 480
rect 454052 354 454080 174558
rect 455420 167952 455472 167958
rect 455420 167894 455472 167900
rect 455432 16574 455460 167894
rect 455432 16546 455736 16574
rect 455708 480 455736 16546
rect 456812 3346 456840 324906
rect 459560 177744 459612 177750
rect 459560 177686 459612 177692
rect 456892 172236 456944 172242
rect 456892 172178 456944 172184
rect 456904 3534 456932 172178
rect 458180 167884 458232 167890
rect 458180 167826 458232 167832
rect 458192 16574 458220 167826
rect 459572 16574 459600 177686
rect 462320 169176 462372 169182
rect 462320 169118 462372 169124
rect 460940 167816 460992 167822
rect 460940 167758 460992 167764
rect 460952 16574 460980 167758
rect 458192 16546 459232 16574
rect 459572 16546 459968 16574
rect 460952 16546 461624 16574
rect 456892 3528 456944 3534
rect 456892 3470 456944 3476
rect 458088 3528 458140 3534
rect 458088 3470 458140 3476
rect 456812 3318 456932 3346
rect 456904 480 456932 3318
rect 458100 480 458128 3470
rect 459204 480 459232 16546
rect 454470 354 454582 480
rect 454052 326 454582 354
rect 454470 -960 454582 326
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 459940 354 459968 16546
rect 461596 480 461624 16546
rect 460358 354 460470 480
rect 459940 326 460470 354
rect 460358 -960 460470 326
rect 461554 -960 461666 480
rect 462332 354 462360 169118
rect 463712 16574 463740 333231
rect 463712 16546 464016 16574
rect 463988 480 464016 16546
rect 465092 3534 465120 338098
rect 474738 336424 474794 336433
rect 474738 336359 474794 336368
rect 467840 336252 467892 336258
rect 467840 336194 467892 336200
rect 465172 159588 465224 159594
rect 465172 159530 465224 159536
rect 465080 3528 465132 3534
rect 465080 3470 465132 3476
rect 465184 480 465212 159530
rect 467852 16574 467880 336194
rect 471980 184204 472032 184210
rect 471980 184146 472032 184152
rect 469220 169108 469272 169114
rect 469220 169050 469272 169056
rect 469232 16574 469260 169050
rect 470600 159520 470652 159526
rect 470600 159462 470652 159468
rect 467852 16546 468248 16574
rect 469232 16546 469904 16574
rect 465908 3528 465960 3534
rect 465908 3470 465960 3476
rect 462750 354 462862 480
rect 462332 326 462862 354
rect 462750 -960 462862 326
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 465920 354 465948 3470
rect 467470 3360 467526 3369
rect 467470 3295 467526 3304
rect 467484 480 467512 3295
rect 466246 354 466358 480
rect 465920 326 466358 354
rect 466246 -960 466358 326
rect 467442 -960 467554 480
rect 468220 354 468248 16546
rect 469876 480 469904 16546
rect 468638 354 468750 480
rect 468220 326 468750 354
rect 468638 -960 468750 326
rect 469834 -960 469946 480
rect 470612 354 470640 159462
rect 471992 16574 472020 184146
rect 473360 170468 473412 170474
rect 473360 170410 473412 170416
rect 471992 16546 472296 16574
rect 472268 480 472296 16546
rect 473372 6914 473400 170410
rect 473452 156800 473504 156806
rect 473452 156742 473504 156748
rect 473464 16574 473492 156742
rect 474752 16574 474780 336359
rect 480258 336288 480314 336297
rect 480258 336223 480314 336232
rect 476120 170400 476172 170406
rect 476120 170342 476172 170348
rect 476132 16574 476160 170342
rect 478880 167748 478932 167754
rect 478880 167690 478932 167696
rect 477500 160948 477552 160954
rect 477500 160890 477552 160896
rect 477512 16574 477540 160890
rect 473464 16546 474136 16574
rect 474752 16546 475792 16574
rect 476132 16546 476528 16574
rect 477512 16546 478184 16574
rect 473372 6886 473492 6914
rect 473464 480 473492 6886
rect 471030 354 471142 480
rect 470612 326 471142 354
rect 471030 -960 471142 326
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474108 354 474136 16546
rect 475764 480 475792 16546
rect 474526 354 474638 480
rect 474108 326 474638 354
rect 474526 -960 474638 326
rect 475722 -960 475834 480
rect 476500 354 476528 16546
rect 478156 480 478184 16546
rect 476918 354 477030 480
rect 476500 326 477030 354
rect 476918 -960 477030 326
rect 478114 -960 478226 480
rect 478892 354 478920 167690
rect 480272 16574 480300 336223
rect 483020 336184 483072 336190
rect 483020 336126 483072 336132
rect 487158 336152 487214 336161
rect 481638 170368 481694 170377
rect 481638 170303 481694 170312
rect 480272 16546 480576 16574
rect 480548 480 480576 16546
rect 481652 6914 481680 170303
rect 481730 160848 481786 160857
rect 481730 160783 481786 160792
rect 481744 16574 481772 160783
rect 483032 16574 483060 336126
rect 487158 336087 487214 336096
rect 500960 336116 501012 336122
rect 484400 172168 484452 172174
rect 484400 172110 484452 172116
rect 484412 16574 484440 172110
rect 485780 169040 485832 169046
rect 485780 168982 485832 168988
rect 485792 16574 485820 168982
rect 481744 16546 482416 16574
rect 483032 16546 484072 16574
rect 484412 16546 484808 16574
rect 485792 16546 486464 16574
rect 481652 6886 481772 6914
rect 481744 480 481772 6886
rect 479310 354 479422 480
rect 478892 326 479422 354
rect 479310 -960 479422 326
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482388 354 482416 16546
rect 484044 480 484072 16546
rect 482806 354 482918 480
rect 482388 326 482918 354
rect 482806 -960 482918 326
rect 484002 -960 484114 480
rect 484780 354 484808 16546
rect 486436 480 486464 16546
rect 485198 354 485310 480
rect 484780 326 485310 354
rect 485198 -960 485310 326
rect 486394 -960 486506 480
rect 487172 354 487200 336087
rect 500960 336058 501012 336064
rect 491300 335096 491352 335102
rect 491300 335038 491352 335044
rect 489920 329180 489972 329186
rect 489920 329122 489972 329128
rect 488540 172100 488592 172106
rect 488540 172042 488592 172048
rect 488552 16574 488580 172042
rect 488552 16546 488856 16574
rect 488828 480 488856 16546
rect 489932 3534 489960 329122
rect 490012 172032 490064 172038
rect 490012 171974 490064 171980
rect 489920 3528 489972 3534
rect 489920 3470 489972 3476
rect 490024 3346 490052 171974
rect 491312 16574 491340 335038
rect 498198 330576 498254 330585
rect 498198 330511 498254 330520
rect 496818 173496 496874 173505
rect 496818 173431 496874 173440
rect 492680 171964 492732 171970
rect 492680 171906 492732 171912
rect 492692 16574 492720 171906
rect 495440 156732 495492 156738
rect 495440 156674 495492 156680
rect 494058 155272 494114 155281
rect 494058 155207 494114 155216
rect 494072 16574 494100 155207
rect 491312 16546 492352 16574
rect 492692 16546 493088 16574
rect 494072 16546 494744 16574
rect 490748 3528 490800 3534
rect 490748 3470 490800 3476
rect 489932 3318 490052 3346
rect 489932 480 489960 3318
rect 487590 354 487702 480
rect 487172 326 487702 354
rect 487590 -960 487702 326
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 490760 354 490788 3470
rect 492324 480 492352 16546
rect 491086 354 491198 480
rect 490760 326 491198 354
rect 491086 -960 491198 326
rect 492282 -960 492394 480
rect 493060 354 493088 16546
rect 494716 480 494744 16546
rect 493478 354 493590 480
rect 493060 326 493590 354
rect 493478 -960 493590 326
rect 494674 -960 494786 480
rect 495452 354 495480 156674
rect 496832 16574 496860 173431
rect 496832 16546 497136 16574
rect 497108 480 497136 16546
rect 498212 3534 498240 330511
rect 499578 174584 499634 174593
rect 499578 174519 499634 174528
rect 498290 156632 498346 156641
rect 498290 156567 498346 156576
rect 498200 3528 498252 3534
rect 498200 3470 498252 3476
rect 498304 3346 498332 156567
rect 499592 16574 499620 174519
rect 500972 16574 501000 336058
rect 518898 336016 518954 336025
rect 518898 335951 518954 335960
rect 509240 335028 509292 335034
rect 509240 334970 509292 334976
rect 503720 177676 503772 177682
rect 503720 177618 503772 177624
rect 502340 156664 502392 156670
rect 502340 156606 502392 156612
rect 502352 16574 502380 156606
rect 499592 16546 500632 16574
rect 500972 16546 501368 16574
rect 502352 16546 503024 16574
rect 499028 3528 499080 3534
rect 499028 3470 499080 3476
rect 498212 3318 498332 3346
rect 498212 480 498240 3318
rect 495870 354 495982 480
rect 495452 326 495982 354
rect 495870 -960 495982 326
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499040 354 499068 3470
rect 500604 480 500632 16546
rect 499366 354 499478 480
rect 499040 326 499478 354
rect 499366 -960 499478 326
rect 500562 -960 500674 480
rect 501340 354 501368 16546
rect 502996 480 503024 16546
rect 501758 354 501870 480
rect 501340 326 501870 354
rect 501758 -960 501870 326
rect 502954 -960 503066 480
rect 503732 354 503760 177618
rect 506480 171896 506532 171902
rect 506480 171838 506532 171844
rect 505100 158024 505152 158030
rect 505100 157966 505152 157972
rect 505112 16574 505140 157966
rect 505112 16546 505416 16574
rect 505388 480 505416 16546
rect 506492 480 506520 171838
rect 506572 162240 506624 162246
rect 506572 162182 506624 162188
rect 506584 16574 506612 162182
rect 507858 157992 507914 158001
rect 507858 157927 507914 157936
rect 507872 16574 507900 157927
rect 509252 16574 509280 334970
rect 516138 334792 516194 334801
rect 516138 334727 516194 334736
rect 514758 327720 514814 327729
rect 514758 327655 514814 327664
rect 512000 326596 512052 326602
rect 512000 326538 512052 326544
rect 510620 177608 510672 177614
rect 510620 177550 510672 177556
rect 510632 16574 510660 177550
rect 506584 16546 507256 16574
rect 507872 16546 508912 16574
rect 509252 16546 509648 16574
rect 510632 16546 511304 16574
rect 504150 354 504262 480
rect 503732 326 504262 354
rect 504150 -960 504262 326
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507228 354 507256 16546
rect 508884 480 508912 16546
rect 507646 354 507758 480
rect 507228 326 507758 354
rect 507646 -960 507758 326
rect 508842 -960 508954 480
rect 509620 354 509648 16546
rect 511276 480 511304 16546
rect 510038 354 510150 480
rect 509620 326 510150 354
rect 510038 -960 510150 326
rect 511234 -960 511346 480
rect 512012 354 512040 326538
rect 513380 171828 513432 171834
rect 513380 171770 513432 171776
rect 512430 354 512542 480
rect 512012 326 512542 354
rect 513392 354 513420 171770
rect 514772 3534 514800 327655
rect 514850 162344 514906 162353
rect 514850 162279 514906 162288
rect 514760 3528 514812 3534
rect 514760 3470 514812 3476
rect 514864 3346 514892 162279
rect 516152 16574 516180 334727
rect 517518 330440 517574 330449
rect 517518 330375 517574 330384
rect 517532 16574 517560 330375
rect 518912 16574 518940 335951
rect 523040 334960 523092 334966
rect 523040 334902 523092 334908
rect 521660 177540 521712 177546
rect 521660 177482 521712 177488
rect 520280 173460 520332 173466
rect 520280 173402 520332 173408
rect 516152 16546 517192 16574
rect 517532 16546 517928 16574
rect 518912 16546 519584 16574
rect 515588 3528 515640 3534
rect 515588 3470 515640 3476
rect 514772 3318 514892 3346
rect 514772 480 514800 3318
rect 513534 354 513646 480
rect 513392 326 513646 354
rect 512430 -960 512542 326
rect 513534 -960 513646 326
rect 514730 -960 514842 480
rect 515600 354 515628 3470
rect 517164 480 517192 16546
rect 515926 354 516038 480
rect 515600 326 516038 354
rect 515926 -960 516038 326
rect 517122 -960 517234 480
rect 517900 354 517928 16546
rect 519556 480 519584 16546
rect 518318 354 518430 480
rect 517900 326 518430 354
rect 518318 -960 518430 326
rect 519514 -960 519626 480
rect 520292 354 520320 173402
rect 520710 354 520822 480
rect 520292 326 520822 354
rect 521672 354 521700 177482
rect 523052 3534 523080 334902
rect 523132 326528 523184 326534
rect 523132 326470 523184 326476
rect 523040 3528 523092 3534
rect 523040 3470 523092 3476
rect 523144 3346 523172 326470
rect 523696 320890 523724 384095
rect 577596 383240 577648 383246
rect 577596 383182 577648 383188
rect 577502 380216 577558 380225
rect 577502 380151 577558 380160
rect 557540 336796 557592 336802
rect 557540 336738 557592 336744
rect 536840 336048 536892 336054
rect 536840 335990 536892 335996
rect 531320 334892 531372 334898
rect 531320 334834 531372 334840
rect 528560 326460 528612 326466
rect 528560 326402 528612 326408
rect 523684 320884 523736 320890
rect 523684 320826 523736 320832
rect 524420 177472 524472 177478
rect 524420 177414 524472 177420
rect 524432 16574 524460 177414
rect 527180 173392 527232 173398
rect 527180 173334 527232 173340
rect 525800 159452 525852 159458
rect 525800 159394 525852 159400
rect 525812 16574 525840 159394
rect 527192 16574 527220 173334
rect 524432 16546 525472 16574
rect 525812 16546 526208 16574
rect 527192 16546 527864 16574
rect 523868 3528 523920 3534
rect 523868 3470 523920 3476
rect 523052 3318 523172 3346
rect 523052 480 523080 3318
rect 521814 354 521926 480
rect 521672 326 521926 354
rect 520710 -960 520822 326
rect 521814 -960 521926 326
rect 523010 -960 523122 480
rect 523880 354 523908 3470
rect 525444 480 525472 16546
rect 524206 354 524318 480
rect 523880 326 524318 354
rect 524206 -960 524318 326
rect 525402 -960 525514 480
rect 526180 354 526208 16546
rect 527836 480 527864 16546
rect 526598 354 526710 480
rect 526180 326 526710 354
rect 526598 -960 526710 326
rect 527794 -960 527906 480
rect 528572 354 528600 326402
rect 529940 159384 529992 159390
rect 529940 159326 529992 159332
rect 528990 354 529102 480
rect 528572 326 529102 354
rect 529952 354 529980 159326
rect 531332 480 531360 334834
rect 535458 332072 535514 332081
rect 535458 332007 535514 332016
rect 534078 173360 534134 173369
rect 534078 173295 534134 173304
rect 531410 162208 531466 162217
rect 531410 162143 531466 162152
rect 531424 16574 531452 162143
rect 532698 159488 532754 159497
rect 532698 159423 532754 159432
rect 532712 16574 532740 159423
rect 534092 16574 534120 173295
rect 535472 16574 535500 332007
rect 536852 16574 536880 335990
rect 538220 334824 538272 334830
rect 538220 334766 538272 334772
rect 531424 16546 532096 16574
rect 532712 16546 533752 16574
rect 534092 16546 534488 16574
rect 535472 16546 536144 16574
rect 536852 16546 537248 16574
rect 530094 354 530206 480
rect 529952 326 530206 354
rect 528990 -960 529102 326
rect 530094 -960 530206 326
rect 531290 -960 531402 480
rect 532068 354 532096 16546
rect 533724 480 533752 16546
rect 532486 354 532598 480
rect 532068 326 532598 354
rect 532486 -960 532598 326
rect 533682 -960 533794 480
rect 534460 354 534488 16546
rect 536116 480 536144 16546
rect 537220 480 537248 16546
rect 534878 354 534990 480
rect 534460 326 534990 354
rect 534878 -960 534990 326
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538232 354 538260 334766
rect 545120 334756 545172 334762
rect 545120 334698 545172 334704
rect 539600 329112 539652 329118
rect 539600 329054 539652 329060
rect 539612 3534 539640 329054
rect 542360 177404 542412 177410
rect 542360 177346 542412 177352
rect 539692 174548 539744 174554
rect 539692 174490 539744 174496
rect 539600 3528 539652 3534
rect 539600 3470 539652 3476
rect 539704 3346 539732 174490
rect 540980 173324 541032 173330
rect 540980 173266 541032 173272
rect 540992 16574 541020 173266
rect 542372 16574 542400 177346
rect 543740 160880 543792 160886
rect 543740 160822 543792 160828
rect 543752 16574 543780 160822
rect 545132 16574 545160 334698
rect 556160 334688 556212 334694
rect 552018 334656 552074 334665
rect 556160 334630 556212 334636
rect 552018 334591 552074 334600
rect 549258 331936 549314 331945
rect 549258 331871 549314 331880
rect 547880 193860 547932 193866
rect 547880 193802 547932 193808
rect 546500 177336 546552 177342
rect 546500 177278 546552 177284
rect 540992 16546 542032 16574
rect 542372 16546 542768 16574
rect 543752 16546 544424 16574
rect 545132 16546 545528 16574
rect 540428 3528 540480 3534
rect 540428 3470 540480 3476
rect 539612 3318 539732 3346
rect 539612 480 539640 3318
rect 538374 354 538486 480
rect 538232 326 538486 354
rect 538374 -960 538486 326
rect 539570 -960 539682 480
rect 540440 354 540468 3470
rect 542004 480 542032 16546
rect 540766 354 540878 480
rect 540440 326 540878 354
rect 540766 -960 540878 326
rect 541962 -960 542074 480
rect 542740 354 542768 16546
rect 544396 480 544424 16546
rect 545500 480 545528 16546
rect 543158 354 543270 480
rect 542740 326 543270 354
rect 543158 -960 543270 326
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546512 354 546540 177278
rect 547892 3534 547920 193802
rect 547972 160812 548024 160818
rect 547972 160754 548024 160760
rect 547880 3528 547932 3534
rect 547880 3470 547932 3476
rect 547984 3346 548012 160754
rect 549272 16574 549300 331871
rect 550638 160712 550694 160721
rect 550638 160647 550694 160656
rect 550652 16574 550680 160647
rect 552032 16574 552060 334591
rect 553398 177304 553454 177313
rect 553398 177239 553454 177248
rect 553412 16574 553440 177239
rect 554780 166320 554832 166326
rect 554780 166262 554832 166268
rect 549272 16546 550312 16574
rect 550652 16546 551048 16574
rect 552032 16546 552704 16574
rect 553412 16546 553808 16574
rect 548708 3528 548760 3534
rect 548708 3470 548760 3476
rect 547892 3318 548012 3346
rect 547892 480 547920 3318
rect 546654 354 546766 480
rect 546512 326 546766 354
rect 546654 -960 546766 326
rect 547850 -960 547962 480
rect 548720 354 548748 3470
rect 550284 480 550312 16546
rect 549046 354 549158 480
rect 548720 326 549158 354
rect 549046 -960 549158 326
rect 550242 -960 550354 480
rect 551020 354 551048 16546
rect 552676 480 552704 16546
rect 553780 480 553808 16546
rect 551438 354 551550 480
rect 551020 326 551550 354
rect 551438 -960 551550 326
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554792 354 554820 166262
rect 556172 480 556200 334630
rect 556252 331968 556304 331974
rect 556252 331910 556304 331916
rect 556264 16574 556292 331910
rect 557552 16574 557580 336738
rect 565820 334620 565872 334626
rect 565820 334562 565872 334568
rect 564440 331900 564492 331906
rect 564440 331842 564492 331848
rect 560300 178900 560352 178906
rect 560300 178842 560352 178848
rect 558920 163532 558972 163538
rect 558920 163474 558972 163480
rect 558932 16574 558960 163474
rect 560312 16574 560340 178842
rect 563060 173256 563112 173262
rect 563060 173198 563112 173204
rect 561680 160744 561732 160750
rect 561680 160686 561732 160692
rect 561692 16574 561720 160686
rect 556264 16546 556936 16574
rect 557552 16546 558592 16574
rect 558932 16546 559328 16574
rect 560312 16546 560432 16574
rect 561692 16546 562088 16574
rect 554934 354 555046 480
rect 554792 326 555046 354
rect 554934 -960 555046 326
rect 556130 -960 556242 480
rect 556908 354 556936 16546
rect 558564 480 558592 16546
rect 557326 354 557438 480
rect 556908 326 557438 354
rect 557326 -960 557438 326
rect 558522 -960 558634 480
rect 559300 354 559328 16546
rect 559718 354 559830 480
rect 559300 326 559830 354
rect 560404 354 560432 16546
rect 562060 480 562088 16546
rect 560822 354 560934 480
rect 560404 326 560934 354
rect 559718 -960 559830 326
rect 560822 -960 560934 326
rect 562018 -960 562130 480
rect 563072 354 563100 173198
rect 564452 480 564480 331842
rect 564532 162172 564584 162178
rect 564532 162114 564584 162120
rect 564544 16574 564572 162114
rect 565832 16574 565860 334562
rect 571338 331800 571394 331809
rect 571338 331735 571394 331744
rect 567200 178832 567252 178838
rect 567200 178774 567252 178780
rect 567212 16574 567240 178774
rect 569958 173224 570014 173233
rect 569958 173159 570014 173168
rect 568578 162072 568634 162081
rect 568578 162007 568634 162016
rect 568592 16574 568620 162007
rect 569972 16574 570000 173159
rect 564544 16546 565216 16574
rect 565832 16546 566872 16574
rect 567212 16546 567608 16574
rect 568592 16546 568712 16574
rect 569972 16546 570368 16574
rect 563214 354 563326 480
rect 563072 326 563326 354
rect 563214 -960 563326 326
rect 564410 -960 564522 480
rect 565188 354 565216 16546
rect 566844 480 566872 16546
rect 565606 354 565718 480
rect 565188 326 565718 354
rect 565606 -960 565718 326
rect 566802 -960 566914 480
rect 567580 354 567608 16546
rect 567998 354 568110 480
rect 567580 326 568110 354
rect 568684 354 568712 16546
rect 570340 480 570368 16546
rect 569102 354 569214 480
rect 568684 326 569214 354
rect 567998 -960 568110 326
rect 569102 -960 569214 326
rect 570298 -960 570410 480
rect 571352 354 571380 331735
rect 572720 330540 572772 330546
rect 572720 330482 572772 330488
rect 572732 480 572760 330482
rect 575480 327752 575532 327758
rect 575480 327694 575532 327700
rect 572812 326392 572864 326398
rect 572812 326334 572864 326340
rect 572824 16574 572852 326334
rect 574100 178764 574152 178770
rect 574100 178706 574152 178712
rect 574112 16574 574140 178706
rect 575492 16574 575520 327694
rect 576860 173188 576912 173194
rect 576860 173130 576912 173136
rect 576872 16574 576900 173130
rect 577516 20670 577544 380151
rect 577608 100706 577636 383182
rect 577686 383072 577742 383081
rect 577686 383007 577742 383016
rect 577700 139398 577728 383007
rect 577792 219230 577820 385018
rect 577870 383208 577926 383217
rect 577870 383143 577926 383152
rect 577780 219224 577832 219230
rect 577780 219166 577832 219172
rect 577884 179382 577912 383143
rect 577976 259418 578004 385086
rect 579988 384600 580040 384606
rect 579988 384542 580040 384548
rect 578056 383172 578108 383178
rect 578056 383114 578108 383120
rect 578068 273222 578096 383114
rect 579896 381608 579948 381614
rect 579896 381550 579948 381556
rect 578146 380352 578202 380361
rect 578146 380287 578202 380296
rect 578160 313274 578188 380287
rect 579908 373994 579936 381550
rect 580000 378826 580028 384542
rect 580540 384532 580592 384538
rect 580540 384474 580592 384480
rect 580446 384024 580502 384033
rect 580446 383959 580502 383968
rect 580264 383104 580316 383110
rect 580264 383046 580316 383052
rect 580080 381540 580132 381546
rect 580080 381482 580132 381488
rect 579988 378820 580040 378826
rect 579988 378762 580040 378768
rect 580092 378298 580120 381482
rect 580172 379500 580224 379506
rect 580172 379442 580224 379448
rect 580184 378457 580212 379442
rect 580170 378448 580226 378457
rect 580170 378383 580226 378392
rect 580092 378270 580212 378298
rect 579908 373966 580120 373994
rect 580092 365129 580120 373966
rect 580078 365120 580134 365129
rect 580078 365055 580134 365064
rect 579988 353252 580040 353258
rect 579988 353194 580040 353200
rect 580000 351937 580028 353194
rect 579986 351928 580042 351937
rect 579986 351863 580042 351872
rect 578148 313268 578200 313274
rect 578148 313210 578200 313216
rect 580080 313268 580132 313274
rect 580080 313210 580132 313216
rect 580092 312089 580120 313210
rect 580078 312080 580134 312089
rect 580078 312015 580134 312024
rect 580184 298761 580212 378270
rect 580276 325281 580304 383046
rect 580354 381032 580410 381041
rect 580354 380967 580410 380976
rect 580262 325272 580318 325281
rect 580262 325207 580318 325216
rect 580264 320884 580316 320890
rect 580264 320826 580316 320832
rect 580170 298752 580226 298761
rect 580170 298687 580226 298696
rect 578056 273216 578108 273222
rect 578056 273158 578108 273164
rect 580080 273216 580132 273222
rect 580080 273158 580132 273164
rect 580092 272241 580120 273158
rect 580078 272232 580134 272241
rect 580078 272167 580134 272176
rect 577964 259412 578016 259418
rect 577964 259354 578016 259360
rect 580080 259412 580132 259418
rect 580080 259354 580132 259360
rect 580092 258913 580120 259354
rect 580078 258904 580134 258913
rect 580078 258839 580134 258848
rect 579712 219224 579764 219230
rect 579712 219166 579764 219172
rect 579724 219065 579752 219166
rect 579710 219056 579766 219065
rect 579710 218991 579766 219000
rect 577872 179376 577924 179382
rect 577872 179318 577924 179324
rect 579712 179376 579764 179382
rect 579712 179318 579764 179324
rect 579724 179217 579752 179318
rect 579710 179208 579766 179217
rect 579710 179143 579766 179152
rect 578240 178696 578292 178702
rect 578240 178638 578292 178644
rect 577688 139392 577740 139398
rect 577688 139334 577740 139340
rect 577596 100700 577648 100706
rect 577596 100642 577648 100648
rect 577504 20664 577556 20670
rect 577504 20606 577556 20612
rect 578252 16574 578280 178638
rect 580172 167000 580224 167006
rect 580172 166942 580224 166948
rect 580184 165889 580212 166942
rect 580170 165880 580226 165889
rect 580170 165815 580226 165824
rect 579620 139392 579672 139398
rect 579618 139360 579620 139369
rect 579672 139360 579674 139369
rect 579618 139295 579674 139304
rect 579712 126948 579764 126954
rect 579712 126890 579764 126896
rect 579724 126041 579752 126890
rect 579710 126032 579766 126041
rect 579710 125967 579766 125976
rect 579620 100700 579672 100706
rect 579620 100642 579672 100648
rect 579632 99521 579660 100642
rect 579618 99512 579674 99521
rect 579618 99447 579674 99456
rect 580276 46345 580304 320826
rect 580368 73001 580396 380967
rect 580460 112849 580488 383959
rect 580552 192545 580580 384474
rect 580630 383888 580686 383897
rect 580630 383823 580686 383832
rect 580538 192536 580594 192545
rect 580538 192471 580594 192480
rect 580538 159352 580594 159361
rect 580538 159287 580594 159296
rect 580446 112840 580502 112849
rect 580446 112775 580502 112784
rect 580552 86193 580580 159287
rect 580644 152697 580672 383823
rect 580724 380996 580776 381002
rect 580724 380938 580776 380944
rect 580736 205737 580764 380938
rect 580908 380928 580960 380934
rect 580908 380870 580960 380876
rect 580816 378820 580868 378826
rect 580816 378762 580868 378768
rect 580828 232393 580856 378762
rect 580920 245585 580948 380870
rect 580906 245576 580962 245585
rect 580906 245511 580962 245520
rect 580814 232384 580870 232393
rect 580814 232319 580870 232328
rect 580722 205728 580778 205737
rect 580722 205663 580778 205672
rect 581000 180124 581052 180130
rect 581000 180066 581052 180072
rect 580630 152688 580686 152697
rect 580630 152623 580686 152632
rect 580538 86184 580594 86193
rect 580538 86119 580594 86128
rect 580354 72992 580410 73001
rect 580354 72927 580410 72936
rect 580262 46336 580318 46345
rect 580262 46271 580318 46280
rect 579712 20664 579764 20670
rect 579712 20606 579764 20612
rect 579724 19825 579752 20606
rect 579710 19816 579766 19825
rect 579710 19751 579766 19760
rect 572824 16546 573496 16574
rect 574112 16546 575152 16574
rect 575492 16546 575888 16574
rect 576872 16546 576992 16574
rect 578252 16546 578648 16574
rect 571494 354 571606 480
rect 571352 326 571606 354
rect 571494 -960 571606 326
rect 572690 -960 572802 480
rect 573468 354 573496 16546
rect 575124 480 575152 16546
rect 573886 354 573998 480
rect 573468 326 573998 354
rect 573886 -960 573998 326
rect 575082 -960 575194 480
rect 575860 354 575888 16546
rect 576278 354 576390 480
rect 575860 326 576390 354
rect 576964 354 576992 16546
rect 578620 480 578648 16546
rect 580172 6860 580224 6866
rect 580172 6802 580224 6808
rect 580184 6633 580212 6802
rect 580170 6624 580226 6633
rect 580170 6559 580226 6568
rect 581012 3534 581040 180066
rect 582380 167680 582432 167686
rect 582380 167622 582432 167628
rect 581092 163600 581144 163606
rect 581092 163542 581144 163548
rect 581000 3528 581052 3534
rect 581000 3470 581052 3476
rect 579804 3460 579856 3466
rect 579804 3402 579856 3408
rect 579816 480 579844 3402
rect 581104 3346 581132 163542
rect 582392 16574 582420 167622
rect 582392 16546 583432 16574
rect 581828 3528 581880 3534
rect 581828 3470 581880 3476
rect 581012 3318 581132 3346
rect 581012 480 581040 3318
rect 577382 354 577494 480
rect 576964 326 577494 354
rect 576278 -960 576390 326
rect 577382 -960 577494 326
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 581840 354 581868 3470
rect 583404 480 583432 16546
rect 582166 354 582278 480
rect 581840 326 582278 354
rect 582166 -960 582278 326
rect 583362 -960 583474 480
<< via2 >>
rect 3422 684256 3478 684312
rect 3422 671200 3478 671256
rect 3422 658144 3478 658200
rect 3422 632068 3424 632088
rect 3424 632068 3476 632088
rect 3476 632068 3478 632088
rect 3422 632032 3478 632068
rect 2778 619132 2834 619168
rect 2778 619112 2780 619132
rect 2780 619112 2832 619132
rect 2832 619112 2834 619132
rect 3238 606056 3294 606112
rect 3422 579944 3478 580000
rect 2778 566888 2834 566944
rect 2778 553832 2834 553888
rect 3330 501744 3386 501800
rect 3330 475632 3386 475688
rect 3330 462576 3386 462632
rect 3330 449520 3386 449576
rect 3146 423544 3202 423600
rect 3146 410488 3202 410544
rect 3330 397468 3332 397488
rect 3332 397468 3384 397488
rect 3384 397468 3386 397488
rect 3330 397432 3386 397468
rect 3514 527856 3570 527912
rect 3606 514800 3662 514856
rect 4802 393896 4858 393952
rect 97814 536968 97870 537024
rect 97630 510176 97686 510232
rect 97538 508272 97594 508328
rect 97722 508544 97778 508600
rect 97906 535880 97962 535936
rect 99194 534248 99250 534304
rect 99102 533160 99158 533216
rect 99010 530168 99066 530224
rect 98918 528536 98974 528592
rect 99286 531528 99342 531584
rect 114466 498072 114522 498128
rect 119342 498072 119398 498128
rect 123390 498092 123446 498128
rect 123390 498072 123392 498092
rect 123392 498072 123444 498092
rect 123444 498072 123446 498092
rect 113086 496848 113142 496904
rect 125230 498072 125286 498128
rect 126794 498072 126850 498128
rect 151726 498072 151782 498128
rect 121366 497392 121422 497448
rect 115478 496868 115534 496904
rect 115478 496848 115480 496868
rect 115480 496848 115532 496868
rect 115532 496848 115534 496868
rect 118606 496848 118662 496904
rect 121274 496848 121330 496904
rect 122746 496848 122802 496904
rect 125506 496848 125562 496904
rect 131026 496848 131082 496904
rect 136546 496848 136602 496904
rect 140686 496848 140742 496904
rect 146206 496848 146262 496904
rect 155866 496848 155922 496904
rect 161386 496848 161442 496904
rect 233790 393896 233846 393952
rect 233790 393372 233846 393408
rect 233790 393352 233792 393372
rect 233792 393352 233844 393372
rect 233844 393352 233846 393372
rect 3146 371320 3202 371376
rect 2962 345344 3018 345400
rect 3146 319232 3202 319288
rect 3330 306176 3386 306232
rect 3238 293120 3294 293176
rect 3330 267144 3386 267200
rect 3330 254088 3386 254144
rect 3330 241032 3386 241088
rect 3330 214920 3386 214976
rect 3330 162832 3386 162888
rect 3330 149776 3386 149832
rect 3054 136720 3110 136776
rect 3330 84632 3386 84688
rect 3330 71576 3386 71632
rect 3330 58520 3386 58576
rect 3514 381112 3570 381168
rect 90362 382608 90418 382664
rect 3790 358400 3846 358456
rect 24858 333240 24914 333296
rect 9678 327664 9734 327720
rect 6918 326304 6974 326360
rect 3698 201864 3754 201920
rect 3606 188808 3662 188864
rect 3606 110608 3662 110664
rect 3514 45464 3570 45520
rect 3514 32408 3570 32464
rect 3514 19352 3570 19408
rect 3422 6432 3478 6488
rect 6458 4800 6514 4856
rect 8758 12960 8814 13016
rect 17038 8880 17094 8936
rect 22558 13096 22614 13152
rect 21822 9016 21878 9072
rect 24214 3304 24270 3360
rect 27618 79328 27674 79384
rect 32402 9152 32458 9208
rect 45558 331744 45614 331800
rect 40222 13232 40278 13288
rect 39578 9288 39634 9344
rect 44270 13368 44326 13424
rect 57978 329024 58034 329080
rect 54942 9424 54998 9480
rect 59358 13504 59414 13560
rect 60830 329160 60886 329216
rect 62118 177248 62174 177304
rect 80058 80688 80114 80744
rect 71502 6160 71558 6216
rect 77390 14456 77446 14512
rect 75918 10240 75974 10296
rect 79230 10376 79286 10432
rect 93858 333376 93914 333432
rect 89166 6296 89222 6352
rect 111798 327936 111854 327992
rect 96618 327800 96674 327856
rect 96250 7520 96306 7576
rect 95146 4936 95202 4992
rect 114558 44784 114614 44840
rect 111614 13640 111670 13696
rect 119894 6432 119950 6488
rect 132498 330384 132554 330440
rect 129738 326440 129794 326496
rect 131762 9560 131818 9616
rect 147678 334600 147734 334656
rect 146298 330520 146354 330576
rect 136454 3440 136510 3496
rect 150438 328072 150494 328128
rect 144734 6568 144790 6624
rect 157798 5072 157854 5128
rect 164238 335960 164294 336016
rect 167182 7656 167238 7712
rect 169574 6704 169630 6760
rect 182822 336368 182878 336424
rect 178866 336232 178922 336288
rect 178682 336096 178738 336152
rect 183558 326576 183614 326632
rect 182914 6840 182970 6896
rect 186318 155352 186374 155408
rect 185030 155216 185086 155272
rect 201498 156576 201554 156632
rect 201590 155488 201646 155544
rect 209870 155624 209926 155680
rect 215298 160656 215354 160712
rect 218150 157936 218206 157992
rect 234066 158344 234122 158400
rect 234342 380432 234398 380488
rect 235262 382744 235318 382800
rect 239218 384376 239274 384432
rect 239678 381928 239734 381984
rect 240782 382064 240838 382120
rect 242162 383832 242218 383888
rect 241426 382336 241482 382392
rect 242438 383016 242494 383072
rect 243266 383152 243322 383208
rect 246026 381928 246082 381984
rect 246302 382064 246358 382120
rect 241886 381656 241942 381712
rect 239954 381384 240010 381440
rect 240506 381384 240562 381440
rect 242714 381384 242770 381440
rect 249062 382336 249118 382392
rect 246302 381520 246358 381576
rect 259642 383560 259698 383616
rect 259642 382880 259698 382936
rect 260194 383560 260250 383616
rect 257894 381792 257950 381848
rect 262126 384240 262182 384296
rect 270866 385056 270922 385112
rect 266450 384104 266506 384160
rect 267646 384412 267648 384432
rect 267648 384412 267700 384432
rect 267700 384412 267702 384432
rect 267646 384376 267702 384412
rect 268198 384376 268254 384432
rect 267554 382744 267610 382800
rect 268658 383968 268714 384024
rect 268382 382608 268438 382664
rect 271418 383288 271474 383344
rect 273074 384648 273130 384704
rect 273442 384784 273498 384840
rect 274546 382064 274602 382120
rect 269210 381792 269266 381848
rect 273902 381792 273958 381848
rect 276754 382472 276810 382528
rect 278042 382608 278098 382664
rect 278410 382336 278466 382392
rect 281078 384512 281134 384568
rect 283976 382064 284032 382120
rect 276110 381792 276166 381848
rect 277766 381792 277822 381848
rect 282458 381792 282514 381848
rect 287886 383696 287942 383752
rect 288530 381928 288586 381984
rect 289358 381928 289414 381984
rect 289726 383968 289782 384024
rect 290002 382064 290058 382120
rect 290922 384104 290978 384160
rect 291106 382744 291162 382800
rect 291842 384412 291844 384432
rect 291844 384412 291896 384432
rect 291896 384412 291898 384432
rect 291842 384376 291898 384412
rect 292118 381928 292174 381984
rect 293912 382064 293968 382120
rect 294878 381928 294934 381984
rect 295614 384920 295670 384976
rect 295338 384820 295340 384840
rect 295340 384820 295392 384840
rect 295392 384820 295394 384840
rect 295338 384784 295394 384820
rect 295706 381928 295762 381984
rect 376942 536968 376998 537024
rect 377034 535880 377090 535936
rect 376942 534248 376998 534304
rect 377034 533160 377090 533216
rect 376942 531528 376998 531584
rect 376942 530168 376998 530224
rect 376850 528572 376852 528592
rect 376852 528572 376904 528592
rect 376904 528572 376906 528592
rect 376850 528536 376906 528572
rect 376942 510176 376998 510232
rect 377034 508544 377090 508600
rect 376758 508272 376814 508328
rect 397458 498072 397514 498128
rect 425058 498072 425114 498128
rect 409878 497664 409934 497720
rect 398930 497256 398986 497312
rect 403162 497256 403218 497312
rect 398838 497140 398894 497176
rect 398838 497120 398840 497140
rect 398840 497120 398892 497140
rect 398892 497120 398894 497140
rect 404358 496984 404414 497040
rect 391938 496848 391994 496904
rect 393318 496848 393374 496904
rect 394698 496848 394754 496904
rect 400218 496848 400274 496904
rect 401598 496848 401654 496904
rect 404450 496848 404506 496904
rect 405738 496848 405794 496904
rect 415398 496848 415454 496904
rect 419538 496848 419594 496904
rect 429198 496848 429254 496904
rect 434718 496848 434774 496904
rect 440238 496848 440294 496904
rect 580170 697176 580226 697232
rect 580170 683848 580226 683904
rect 580170 670692 580172 670712
rect 580172 670692 580224 670712
rect 580224 670692 580226 670712
rect 580170 670656 580226 670692
rect 580170 644000 580226 644056
rect 580170 630808 580226 630864
rect 580170 617480 580226 617536
rect 579802 590960 579858 591016
rect 580354 577632 580410 577688
rect 580262 564304 580318 564360
rect 579618 511264 579674 511320
rect 580170 484608 580226 484664
rect 579986 471416 580042 471472
rect 580170 458088 580226 458144
rect 579618 431568 579674 431624
rect 579710 418240 579766 418296
rect 579986 404912 580042 404968
rect 580446 537784 580502 537840
rect 580538 524456 580594 524512
rect 295982 384920 296038 384976
rect 296258 381928 296314 381984
rect 296626 383696 296682 383752
rect 245474 381384 245530 381440
rect 246026 381384 246082 381440
rect 237378 328208 237434 328264
rect 235998 159296 236054 159352
rect 237470 214548 237472 214568
rect 237472 214548 237524 214568
rect 237524 214548 237526 214568
rect 237470 214512 237526 214548
rect 239586 161064 239642 161120
rect 238758 158072 238814 158128
rect 239862 160792 239918 160848
rect 241150 161336 241206 161392
rect 241242 161200 241298 161256
rect 242530 335416 242586 335472
rect 243542 331880 243598 331936
rect 243818 335688 243874 335744
rect 244646 338272 244702 338328
rect 244370 337864 244426 337920
rect 291014 338136 291070 338192
rect 244646 336096 244702 336152
rect 244738 329024 244794 329080
rect 245428 337898 245484 337954
rect 244922 337592 244978 337648
rect 245014 336368 245070 336424
rect 245796 337898 245852 337954
rect 245980 337898 246036 337954
rect 246164 337898 246220 337954
rect 246118 337728 246174 337784
rect 246532 337898 246588 337954
rect 246992 337864 247048 337920
rect 247452 337864 247508 337920
rect 245750 337456 245806 337512
rect 245566 336640 245622 336696
rect 245106 336232 245162 336288
rect 245474 336096 245530 336152
rect 245014 335824 245070 335880
rect 245382 335552 245438 335608
rect 245566 335688 245622 335744
rect 245474 335416 245530 335472
rect 245934 334736 245990 334792
rect 246946 337728 247002 337784
rect 245566 160520 245622 160576
rect 245750 9016 245806 9072
rect 246854 336096 246910 336152
rect 247038 337592 247094 337648
rect 247222 337748 247278 337784
rect 247222 337728 247224 337748
rect 247224 337728 247276 337748
rect 247276 337728 247278 337748
rect 247130 335280 247186 335336
rect 245842 8880 245898 8936
rect 247314 333240 247370 333296
rect 247912 337898 247968 337954
rect 247406 333104 247462 333160
rect 247958 337728 248014 337784
rect 248556 337864 248612 337920
rect 248694 337728 248750 337784
rect 247866 9288 247922 9344
rect 248510 333240 248566 333296
rect 248326 158208 248382 158264
rect 248234 153720 248290 153776
rect 247958 9152 248014 9208
rect 249568 337898 249624 337954
rect 249936 337864 249992 337920
rect 250212 337764 250214 337784
rect 250214 337764 250266 337784
rect 250266 337764 250268 337784
rect 248970 331744 249026 331800
rect 248602 9424 248658 9480
rect 249430 337592 249486 337648
rect 250212 337728 250268 337764
rect 250396 337898 250452 337954
rect 250948 337898 251004 337954
rect 251224 337898 251280 337954
rect 250258 337592 250314 337648
rect 249522 329160 249578 329216
rect 249982 337456 250038 337512
rect 251592 337864 251648 337920
rect 251960 337898 252016 337954
rect 250810 337456 250866 337512
rect 251086 337320 251142 337376
rect 251454 333376 251510 333432
rect 251270 333240 251326 333296
rect 249890 6160 249946 6216
rect 251914 337728 251970 337784
rect 252420 337898 252476 337954
rect 252282 337728 252338 337784
rect 252880 337864 252936 337920
rect 252788 337728 252844 337784
rect 253064 337864 253120 337920
rect 252650 334736 252706 334792
rect 253202 337728 253258 337784
rect 253202 336640 253258 336696
rect 253984 337898 254040 337954
rect 254168 337898 254224 337954
rect 254352 337898 254408 337954
rect 254996 337898 255052 337954
rect 255456 337898 255512 337954
rect 255640 337898 255696 337954
rect 253938 337340 253994 337376
rect 253938 337320 253940 337340
rect 253940 337320 253992 337340
rect 253992 337320 253994 337340
rect 254122 334464 254178 334520
rect 254214 332832 254270 332888
rect 254398 337456 254454 337512
rect 253110 158616 253166 158672
rect 251730 6296 251786 6352
rect 255548 337762 255604 337818
rect 254490 6840 254546 6896
rect 255824 337864 255880 337920
rect 256100 337864 256156 337920
rect 255594 337592 255650 337648
rect 254766 6432 254822 6488
rect 255870 337456 255926 337512
rect 255962 335824 256018 335880
rect 256744 337898 256800 337954
rect 256560 337830 256616 337886
rect 256514 337592 256570 337648
rect 255686 159432 255742 159488
rect 255226 3304 255282 3360
rect 256054 326304 256110 326360
rect 257480 337864 257536 337920
rect 257756 337864 257812 337920
rect 256790 334600 256846 334656
rect 256146 6568 256202 6624
rect 257066 335280 257122 335336
rect 257618 337728 257674 337784
rect 257342 334736 257398 334792
rect 257526 337592 257582 337648
rect 257618 333920 257674 333976
rect 256698 152360 256754 152416
rect 256698 143520 256754 143576
rect 257894 332152 257950 332208
rect 257342 163376 257398 163432
rect 257250 148280 257306 148336
rect 257250 139440 257306 139496
rect 256790 134680 256846 134736
rect 256790 130600 256846 130656
rect 256790 125840 256846 125896
rect 256790 121760 256846 121816
rect 256790 112920 256846 112976
rect 256790 104080 256846 104136
rect 257434 155896 257490 155952
rect 257618 155080 257674 155136
rect 257802 141888 257858 141944
rect 257802 132504 257858 132560
rect 257802 132368 257858 132424
rect 257802 122848 257858 122904
rect 257802 122712 257858 122768
rect 257802 113192 257858 113248
rect 257802 113056 257858 113112
rect 257802 103536 257858 103592
rect 257802 103400 257858 103456
rect 258308 337864 258364 337920
rect 258216 337728 258272 337784
rect 258354 336504 258410 336560
rect 258262 336096 258318 336152
rect 258078 335960 258134 336016
rect 258170 335824 258226 335880
rect 257802 93880 257858 93936
rect 257986 93744 258042 93800
rect 257986 84224 258042 84280
rect 257986 84088 258042 84144
rect 257986 74568 258042 74624
rect 257986 74432 258042 74488
rect 257986 64912 258042 64968
rect 257986 64776 258042 64832
rect 257986 55256 258042 55312
rect 257986 55120 258042 55176
rect 257986 45600 258042 45656
rect 257986 45464 258042 45520
rect 257986 35944 258042 36000
rect 257986 35808 258042 35864
rect 257986 26288 258042 26344
rect 257986 26152 258042 26208
rect 257986 16632 258042 16688
rect 257986 16496 258042 16552
rect 258446 158752 258502 158808
rect 257986 6976 258042 7032
rect 259320 337898 259376 337954
rect 259780 337898 259836 337954
rect 259274 337728 259330 337784
rect 260148 337864 260204 337920
rect 259872 337764 259874 337784
rect 259874 337764 259926 337784
rect 259926 337764 259928 337784
rect 259872 337728 259928 337764
rect 259550 335688 259606 335744
rect 259642 334464 259698 334520
rect 258998 158480 259054 158536
rect 260102 337592 260158 337648
rect 260976 337864 261032 337920
rect 260286 155660 260288 155680
rect 260288 155660 260340 155680
rect 260340 155660 260342 155680
rect 260286 155624 260342 155660
rect 261528 337898 261584 337954
rect 261206 337592 261262 337648
rect 261022 335280 261078 335336
rect 261482 337456 261538 337512
rect 261390 160656 261446 160712
rect 261988 337898 262044 337954
rect 262356 337728 262412 337784
rect 262632 337898 262688 337954
rect 262816 337864 262872 337920
rect 263184 337898 263240 337954
rect 262126 337592 262182 337648
rect 262310 337592 262366 337648
rect 262586 335824 262642 335880
rect 263046 337728 263102 337784
rect 263920 337864 263976 337920
rect 263736 337728 263792 337784
rect 263874 336640 263930 336696
rect 264472 337864 264528 337920
rect 263506 331064 263562 331120
rect 263506 321544 263562 321600
rect 264702 337728 264758 337784
rect 265116 337898 265172 337954
rect 265392 337864 265448 337920
rect 265576 337898 265632 337954
rect 265438 337728 265494 337784
rect 265070 335416 265126 335472
rect 265254 335552 265310 335608
rect 266128 337830 266184 337886
rect 265530 337592 265586 337648
rect 265438 335416 265494 335472
rect 266082 337456 266138 337512
rect 266680 337864 266736 337920
rect 266358 336776 266414 336832
rect 266542 337592 266598 337648
rect 267600 337864 267656 337920
rect 267462 336640 267518 336696
rect 267968 337864 268024 337920
rect 266450 155624 266506 155680
rect 268014 337728 268070 337784
rect 268704 337864 268760 337920
rect 268750 337728 268806 337784
rect 268842 335552 268898 335608
rect 269026 335688 269082 335744
rect 268934 335416 268990 335472
rect 269026 158616 269082 158672
rect 269486 335416 269542 335472
rect 269578 161336 269634 161392
rect 269670 160792 269726 160848
rect 270452 337864 270508 337920
rect 270406 337764 270408 337784
rect 270408 337764 270460 337784
rect 270460 337764 270462 337784
rect 270406 337728 270462 337764
rect 270820 337898 270876 337954
rect 271280 337728 271336 337784
rect 269854 161200 269910 161256
rect 269762 160520 269818 160576
rect 269302 155760 269358 155816
rect 271142 337456 271198 337512
rect 271694 336232 271750 336288
rect 272384 337864 272440 337920
rect 271786 335416 271842 335472
rect 272476 337728 272532 337784
rect 272430 336096 272486 336152
rect 272338 161064 272394 161120
rect 273672 337864 273728 337920
rect 273166 337592 273222 337648
rect 269394 155352 269450 155408
rect 274408 337898 274464 337954
rect 274592 337864 274648 337920
rect 273810 337592 273866 337648
rect 274270 337456 274326 337512
rect 275236 337898 275292 337954
rect 275696 337864 275752 337920
rect 274822 337592 274878 337648
rect 274638 337456 274694 337512
rect 275420 337728 275476 337784
rect 274638 335280 274694 335336
rect 274454 333240 274510 333296
rect 275006 335280 275062 335336
rect 275650 337456 275706 337512
rect 275834 337592 275890 337648
rect 276432 337728 276488 337784
rect 277076 337898 277132 337954
rect 276478 337592 276534 337648
rect 276570 333648 276626 333704
rect 278272 337898 278328 337954
rect 277122 335960 277178 336016
rect 278226 337728 278282 337784
rect 278548 337898 278604 337954
rect 278824 337864 278880 337920
rect 278640 337728 278696 337784
rect 278410 337592 278466 337648
rect 278410 333512 278466 333568
rect 278502 333240 278558 333296
rect 279928 337864 279984 337920
rect 280112 337830 280168 337886
rect 279974 337764 279976 337784
rect 279976 337764 280028 337784
rect 280028 337764 280030 337784
rect 279974 337728 280030 337764
rect 280388 337864 280444 337920
rect 280848 337898 280904 337954
rect 281492 337864 281548 337920
rect 279882 336252 279938 336288
rect 279882 336232 279884 336252
rect 279884 336232 279936 336252
rect 279936 336232 279938 336252
rect 279790 333376 279846 333432
rect 280342 336640 280398 336696
rect 280710 336268 280712 336288
rect 280712 336268 280764 336288
rect 280764 336268 280766 336288
rect 280710 336232 280766 336268
rect 280894 336776 280950 336832
rect 280894 336640 280950 336696
rect 280802 333240 280858 333296
rect 280986 335688 281042 335744
rect 281354 337592 281410 337648
rect 282044 337864 282100 337920
rect 282320 337864 282376 337920
rect 281998 337728 282054 337784
rect 277398 158344 277454 158400
rect 281906 336776 281962 336832
rect 282780 337864 282836 337920
rect 282918 337456 282974 337512
rect 282734 336232 282790 336288
rect 282458 333784 282514 333840
rect 283194 336640 283250 336696
rect 283884 337864 283940 337920
rect 283470 336776 283526 336832
rect 283470 335416 283526 335472
rect 284436 337864 284492 337920
rect 284022 335824 284078 335880
rect 284298 337592 284354 337648
rect 284206 335552 284262 335608
rect 283930 335416 283986 335472
rect 284114 335416 284170 335472
rect 284988 337728 285044 337784
rect 285632 337864 285688 337920
rect 285310 336776 285366 336832
rect 285816 337728 285872 337784
rect 286184 337864 286240 337920
rect 285586 336368 285642 336424
rect 285494 335552 285550 335608
rect 285310 335416 285366 335472
rect 285862 337456 285918 337512
rect 285770 336096 285826 336152
rect 285218 334736 285274 334792
rect 284390 157936 284446 157992
rect 286138 337456 286194 337512
rect 286920 337898 286976 337954
rect 286736 337728 286792 337784
rect 287288 337864 287344 337920
rect 287472 337898 287528 337954
rect 287748 337898 287804 337954
rect 288116 337898 288172 337954
rect 288392 337898 288448 337954
rect 286874 335144 286930 335200
rect 287334 337728 287390 337784
rect 288208 337764 288210 337784
rect 288210 337764 288262 337784
rect 288262 337764 288264 337784
rect 287426 337592 287482 337648
rect 288208 337728 288264 337764
rect 287610 336368 287666 336424
rect 287610 335960 287666 336016
rect 288530 337456 288586 337512
rect 288254 334600 288310 334656
rect 287702 194520 287758 194576
rect 288944 337898 289000 337954
rect 289128 337728 289184 337784
rect 289588 337898 289644 337954
rect 289772 337898 289828 337954
rect 290140 337898 290196 337954
rect 290416 337898 290472 337954
rect 288898 337592 288954 337648
rect 288714 337184 288770 337240
rect 288714 326712 288770 326768
rect 288714 326440 288770 326496
rect 289726 335008 289782 335064
rect 290094 336640 290150 336696
rect 290094 336096 290150 336152
rect 290278 337728 290334 337784
rect 290646 335416 290702 335472
rect 293958 338000 294014 338056
rect 292670 337864 292726 337920
rect 292854 337184 292910 337240
rect 292670 336640 292726 336696
rect 291198 332016 291254 332072
rect 289634 158344 289690 158400
rect 295982 335416 296038 335472
rect 296626 335280 296682 335336
rect 296626 325760 296682 325816
rect 296626 325624 296682 325680
rect 296626 316104 296682 316160
rect 296626 315968 296682 316024
rect 296626 306448 296682 306504
rect 296626 306312 296682 306368
rect 296626 296792 296682 296848
rect 296626 296656 296682 296712
rect 296626 287136 296682 287192
rect 296626 287000 296682 287056
rect 296626 277480 296682 277536
rect 296626 277344 296682 277400
rect 296626 267824 296682 267880
rect 296626 267688 296682 267744
rect 296626 248376 296682 248432
rect 296626 248240 296682 248296
rect 296626 238720 296682 238776
rect 296626 238584 296682 238640
rect 296626 229064 296682 229120
rect 296626 228928 296682 228984
rect 296626 219408 296682 219464
rect 296626 219272 296682 219328
rect 296626 209752 296682 209808
rect 296626 209616 296682 209672
rect 296626 200096 296682 200152
rect 296626 199960 296682 200016
rect 296626 190440 296682 190496
rect 296626 190304 296682 190360
rect 296626 180784 296682 180840
rect 296626 180648 296682 180704
rect 296626 171128 296682 171184
rect 296626 170992 296682 171048
rect 296626 161472 296682 161528
rect 298006 158616 298062 158672
rect 301042 380568 301098 380624
rect 301134 380432 301190 380488
rect 343730 384376 343786 384432
rect 301778 161336 301834 161392
rect 302514 157800 302570 157856
rect 311162 336640 311218 336696
rect 310886 158480 310942 158536
rect 335358 214512 335414 214568
rect 343638 158344 343694 158400
rect 343730 157392 343786 157448
rect 284022 155624 284078 155680
rect 273166 155352 273222 155408
rect 342810 100680 342866 100736
rect 260010 97552 260066 97608
rect 272246 97688 272302 97744
rect 288990 97824 289046 97880
rect 330850 97824 330906 97880
rect 274822 3848 274878 3904
rect 306746 3712 306802 3768
rect 310242 3576 310298 3632
rect 313830 3440 313886 3496
rect 317326 3304 317382 3360
rect 335082 3304 335138 3360
rect 336278 3032 336334 3088
rect 343362 3848 343418 3904
rect 339866 3712 339922 3768
rect 338670 3576 338726 3632
rect 342166 3304 342222 3360
rect 340970 3168 341026 3224
rect 344098 103400 344154 103456
rect 344190 3984 344246 4040
rect 523682 384104 523738 384160
rect 347042 381656 347098 381712
rect 344650 151680 344706 151736
rect 344650 148280 344706 148336
rect 345110 147600 345166 147656
rect 345018 134000 345074 134056
rect 344926 129784 344982 129840
rect 344466 3576 344522 3632
rect 345018 116320 345074 116376
rect 345386 179968 345442 180024
rect 345294 158208 345350 158264
rect 345202 107480 345258 107536
rect 344834 3576 344890 3632
rect 344558 3440 344614 3496
rect 345478 170448 345534 170504
rect 345570 129920 345626 129976
rect 345478 125160 345534 125216
rect 345386 112240 345442 112296
rect 345846 155488 345902 155544
rect 345754 138760 345810 138816
rect 345294 3440 345350 3496
rect 344834 3168 344890 3224
rect 346490 3304 346546 3360
rect 356702 383696 356758 383752
rect 348330 161200 348386 161256
rect 348146 158072 348202 158128
rect 347134 3032 347190 3088
rect 349434 160928 349490 160984
rect 349434 3576 349490 3632
rect 349894 155624 349950 155680
rect 356058 155352 356114 155408
rect 349710 3712 349766 3768
rect 407762 381248 407818 381304
rect 382922 336504 382978 336560
rect 373998 320728 374054 320784
rect 374090 174664 374146 174720
rect 375378 165008 375434 165064
rect 391938 333648 391994 333704
rect 390558 164872 390614 164928
rect 407210 175888 407266 175944
rect 427818 333512 427874 333568
rect 409878 159568 409934 159624
rect 425058 166504 425114 166560
rect 426438 166368 426494 166424
rect 445758 333376 445814 333432
rect 444378 186904 444434 186960
rect 447138 166232 447194 166288
rect 463698 333240 463754 333296
rect 474738 336368 474794 336424
rect 467470 3304 467526 3360
rect 480258 336232 480314 336288
rect 481638 170312 481694 170368
rect 481730 160792 481786 160848
rect 487158 336096 487214 336152
rect 498198 330520 498254 330576
rect 496818 173440 496874 173496
rect 494058 155216 494114 155272
rect 499578 174528 499634 174584
rect 498290 156576 498346 156632
rect 518898 335960 518954 336016
rect 507858 157936 507914 157992
rect 516138 334736 516194 334792
rect 514758 327664 514814 327720
rect 514850 162288 514906 162344
rect 517518 330384 517574 330440
rect 577502 380160 577558 380216
rect 535458 332016 535514 332072
rect 534078 173304 534134 173360
rect 531410 162152 531466 162208
rect 532698 159432 532754 159488
rect 552018 334600 552074 334656
rect 549258 331880 549314 331936
rect 550638 160656 550694 160712
rect 553398 177248 553454 177304
rect 571338 331744 571394 331800
rect 569958 173168 570014 173224
rect 568578 162016 568634 162072
rect 577686 383016 577742 383072
rect 577870 383152 577926 383208
rect 578146 380296 578202 380352
rect 580446 383968 580502 384024
rect 580170 378392 580226 378448
rect 580078 365064 580134 365120
rect 579986 351872 580042 351928
rect 580078 312024 580134 312080
rect 580354 380976 580410 381032
rect 580262 325216 580318 325272
rect 580170 298696 580226 298752
rect 580078 272176 580134 272232
rect 580078 258848 580134 258904
rect 579710 219000 579766 219056
rect 579710 179152 579766 179208
rect 580170 165824 580226 165880
rect 579618 139340 579620 139360
rect 579620 139340 579672 139360
rect 579672 139340 579674 139360
rect 579618 139304 579674 139340
rect 579710 125976 579766 126032
rect 579618 99456 579674 99512
rect 580630 383832 580686 383888
rect 580538 192480 580594 192536
rect 580538 159296 580594 159352
rect 580446 112784 580502 112840
rect 580906 245520 580962 245576
rect 580814 232328 580870 232384
rect 580722 205672 580778 205728
rect 580630 152632 580686 152688
rect 580538 86128 580594 86184
rect 580354 72936 580410 72992
rect 580262 46280 580318 46336
rect 579710 19760 579766 19816
rect 580170 6568 580226 6624
<< metal3 >>
rect -960 697220 480 697460
rect 580165 697234 580231 697237
rect 583520 697234 584960 697324
rect 580165 697232 584960 697234
rect 580165 697176 580170 697232
rect 580226 697176 584960 697232
rect 580165 697174 584960 697176
rect 580165 697171 580231 697174
rect 583520 697084 584960 697174
rect -960 684314 480 684404
rect 3417 684314 3483 684317
rect -960 684312 3483 684314
rect -960 684256 3422 684312
rect 3478 684256 3483 684312
rect -960 684254 3483 684256
rect -960 684164 480 684254
rect 3417 684251 3483 684254
rect 580165 683906 580231 683909
rect 583520 683906 584960 683996
rect 580165 683904 584960 683906
rect 580165 683848 580170 683904
rect 580226 683848 584960 683904
rect 580165 683846 584960 683848
rect 580165 683843 580231 683846
rect 583520 683756 584960 683846
rect -960 671258 480 671348
rect 3417 671258 3483 671261
rect -960 671256 3483 671258
rect -960 671200 3422 671256
rect 3478 671200 3483 671256
rect -960 671198 3483 671200
rect -960 671108 480 671198
rect 3417 671195 3483 671198
rect 580165 670714 580231 670717
rect 583520 670714 584960 670804
rect 580165 670712 584960 670714
rect 580165 670656 580170 670712
rect 580226 670656 584960 670712
rect 580165 670654 584960 670656
rect 580165 670651 580231 670654
rect 583520 670564 584960 670654
rect -960 658202 480 658292
rect 3417 658202 3483 658205
rect -960 658200 3483 658202
rect -960 658144 3422 658200
rect 3478 658144 3483 658200
rect -960 658142 3483 658144
rect -960 658052 480 658142
rect 3417 658139 3483 658142
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 580165 644058 580231 644061
rect 583520 644058 584960 644148
rect 580165 644056 584960 644058
rect 580165 644000 580170 644056
rect 580226 644000 584960 644056
rect 580165 643998 584960 644000
rect 580165 643995 580231 643998
rect 583520 643908 584960 643998
rect -960 632090 480 632180
rect 3417 632090 3483 632093
rect -960 632088 3483 632090
rect -960 632032 3422 632088
rect 3478 632032 3483 632088
rect -960 632030 3483 632032
rect -960 631940 480 632030
rect 3417 632027 3483 632030
rect 580165 630866 580231 630869
rect 583520 630866 584960 630956
rect 580165 630864 584960 630866
rect 580165 630808 580170 630864
rect 580226 630808 584960 630864
rect 580165 630806 584960 630808
rect 580165 630803 580231 630806
rect 583520 630716 584960 630806
rect -960 619170 480 619260
rect 2773 619170 2839 619173
rect -960 619168 2839 619170
rect -960 619112 2778 619168
rect 2834 619112 2839 619168
rect -960 619110 2839 619112
rect -960 619020 480 619110
rect 2773 619107 2839 619110
rect 580165 617538 580231 617541
rect 583520 617538 584960 617628
rect 580165 617536 584960 617538
rect 580165 617480 580170 617536
rect 580226 617480 584960 617536
rect 580165 617478 584960 617480
rect 580165 617475 580231 617478
rect 583520 617388 584960 617478
rect -960 606114 480 606204
rect 3233 606114 3299 606117
rect -960 606112 3299 606114
rect -960 606056 3238 606112
rect 3294 606056 3299 606112
rect -960 606054 3299 606056
rect -960 605964 480 606054
rect 3233 606051 3299 606054
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 579797 591018 579863 591021
rect 583520 591018 584960 591108
rect 579797 591016 584960 591018
rect 579797 590960 579802 591016
rect 579858 590960 584960 591016
rect 579797 590958 584960 590960
rect 579797 590955 579863 590958
rect 583520 590868 584960 590958
rect -960 580002 480 580092
rect 3417 580002 3483 580005
rect -960 580000 3483 580002
rect -960 579944 3422 580000
rect 3478 579944 3483 580000
rect -960 579942 3483 579944
rect -960 579852 480 579942
rect 3417 579939 3483 579942
rect 580349 577690 580415 577693
rect 583520 577690 584960 577780
rect 580349 577688 584960 577690
rect 580349 577632 580354 577688
rect 580410 577632 584960 577688
rect 580349 577630 584960 577632
rect 580349 577627 580415 577630
rect 583520 577540 584960 577630
rect -960 566946 480 567036
rect 2773 566946 2839 566949
rect -960 566944 2839 566946
rect -960 566888 2778 566944
rect 2834 566888 2839 566944
rect -960 566886 2839 566888
rect -960 566796 480 566886
rect 2773 566883 2839 566886
rect 580257 564362 580323 564365
rect 583520 564362 584960 564452
rect 580257 564360 584960 564362
rect 580257 564304 580262 564360
rect 580318 564304 584960 564360
rect 580257 564302 584960 564304
rect 580257 564299 580323 564302
rect 583520 564212 584960 564302
rect -960 553890 480 553980
rect 2773 553890 2839 553893
rect -960 553888 2839 553890
rect -960 553832 2778 553888
rect 2834 553832 2839 553888
rect -960 553830 2839 553832
rect -960 553740 480 553830
rect 2773 553827 2839 553830
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 580441 537842 580507 537845
rect 583520 537842 584960 537932
rect 580441 537840 584960 537842
rect 580441 537784 580446 537840
rect 580502 537784 584960 537840
rect 580441 537782 584960 537784
rect 580441 537779 580507 537782
rect 583520 537692 584960 537782
rect 97809 537026 97875 537029
rect 99422 537026 100004 537060
rect 97809 537024 100004 537026
rect 97809 536968 97814 537024
rect 97870 537000 100004 537024
rect 376937 537026 377003 537029
rect 379470 537026 380052 537060
rect 376937 537024 380052 537026
rect 97870 536968 99482 537000
rect 97809 536966 99482 536968
rect 376937 536968 376942 537024
rect 376998 537000 380052 537024
rect 376998 536968 379530 537000
rect 376937 536966 379530 536968
rect 97809 536963 97875 536966
rect 376937 536963 377003 536966
rect 97901 535938 97967 535941
rect 99422 535938 100004 535972
rect 97901 535936 100004 535938
rect 97901 535880 97906 535936
rect 97962 535912 100004 535936
rect 377029 535938 377095 535941
rect 379470 535938 380052 535972
rect 377029 535936 380052 535938
rect 97962 535880 99482 535912
rect 97901 535878 99482 535880
rect 377029 535880 377034 535936
rect 377090 535912 380052 535936
rect 377090 535880 379530 535912
rect 377029 535878 379530 535880
rect 97901 535875 97967 535878
rect 377029 535875 377095 535878
rect 99189 534306 99255 534309
rect 99422 534306 100004 534340
rect 99189 534304 100004 534306
rect 99189 534248 99194 534304
rect 99250 534280 100004 534304
rect 376937 534306 377003 534309
rect 379470 534306 380052 534340
rect 376937 534304 380052 534306
rect 99250 534248 99482 534280
rect 99189 534246 99482 534248
rect 376937 534248 376942 534304
rect 376998 534280 380052 534304
rect 376998 534248 379530 534280
rect 376937 534246 379530 534248
rect 99189 534243 99255 534246
rect 376937 534243 377003 534246
rect 99097 533218 99163 533221
rect 99422 533218 100004 533252
rect 99097 533216 100004 533218
rect 99097 533160 99102 533216
rect 99158 533192 100004 533216
rect 377029 533218 377095 533221
rect 379470 533218 380052 533252
rect 377029 533216 380052 533218
rect 99158 533160 99482 533192
rect 99097 533158 99482 533160
rect 377029 533160 377034 533216
rect 377090 533192 380052 533216
rect 377090 533160 379530 533192
rect 377029 533158 379530 533160
rect 99097 533155 99163 533158
rect 377029 533155 377095 533158
rect 99281 531586 99347 531589
rect 99422 531586 100004 531620
rect 99281 531584 100004 531586
rect 99281 531528 99286 531584
rect 99342 531560 100004 531584
rect 376937 531586 377003 531589
rect 379470 531586 380052 531620
rect 376937 531584 380052 531586
rect 99342 531528 99482 531560
rect 99281 531526 99482 531528
rect 376937 531528 376942 531584
rect 376998 531560 380052 531584
rect 376998 531528 379530 531560
rect 376937 531526 379530 531528
rect 99281 531523 99347 531526
rect 376937 531523 377003 531526
rect 99005 530226 99071 530229
rect 99422 530226 100004 530260
rect 99005 530224 100004 530226
rect 99005 530168 99010 530224
rect 99066 530200 100004 530224
rect 376937 530226 377003 530229
rect 379470 530226 380052 530260
rect 376937 530224 380052 530226
rect 99066 530168 99482 530200
rect 99005 530166 99482 530168
rect 376937 530168 376942 530224
rect 376998 530200 380052 530224
rect 376998 530168 379530 530200
rect 376937 530166 379530 530168
rect 99005 530163 99071 530166
rect 376937 530163 377003 530166
rect 98913 528594 98979 528597
rect 99422 528594 100004 528628
rect 98913 528592 100004 528594
rect 98913 528536 98918 528592
rect 98974 528568 100004 528592
rect 376845 528594 376911 528597
rect 379470 528594 380052 528628
rect 376845 528592 380052 528594
rect 98974 528536 99482 528568
rect 98913 528534 99482 528536
rect 376845 528536 376850 528592
rect 376906 528568 380052 528592
rect 376906 528536 379530 528568
rect 376845 528534 379530 528536
rect 98913 528531 98979 528534
rect 376845 528531 376911 528534
rect -960 527914 480 528004
rect 3509 527914 3575 527917
rect -960 527912 3575 527914
rect -960 527856 3514 527912
rect 3570 527856 3575 527912
rect -960 527854 3575 527856
rect -960 527764 480 527854
rect 3509 527851 3575 527854
rect 580533 524514 580599 524517
rect 583520 524514 584960 524604
rect 580533 524512 584960 524514
rect 580533 524456 580538 524512
rect 580594 524456 584960 524512
rect 580533 524454 584960 524456
rect 580533 524451 580599 524454
rect 583520 524364 584960 524454
rect -960 514858 480 514948
rect 3601 514858 3667 514861
rect -960 514856 3667 514858
rect -960 514800 3606 514856
rect 3662 514800 3667 514856
rect -960 514798 3667 514800
rect -960 514708 480 514798
rect 3601 514795 3667 514798
rect 579613 511322 579679 511325
rect 583520 511322 584960 511412
rect 579613 511320 584960 511322
rect 579613 511264 579618 511320
rect 579674 511264 584960 511320
rect 579613 511262 584960 511264
rect 579613 511259 579679 511262
rect 583520 511172 584960 511262
rect 97625 510234 97691 510237
rect 99422 510234 100004 510268
rect 97625 510232 100004 510234
rect 97625 510176 97630 510232
rect 97686 510208 100004 510232
rect 376937 510234 377003 510237
rect 379470 510234 380052 510268
rect 376937 510232 380052 510234
rect 97686 510176 99482 510208
rect 97625 510174 99482 510176
rect 376937 510176 376942 510232
rect 376998 510208 380052 510232
rect 376998 510176 379530 510208
rect 376937 510174 379530 510176
rect 97625 510171 97691 510174
rect 376937 510171 377003 510174
rect 97717 508602 97783 508605
rect 99422 508602 100004 508636
rect 97717 508600 100004 508602
rect 97717 508544 97722 508600
rect 97778 508576 100004 508600
rect 377029 508602 377095 508605
rect 379470 508602 380052 508636
rect 377029 508600 380052 508602
rect 97778 508544 99482 508576
rect 97717 508542 99482 508544
rect 377029 508544 377034 508600
rect 377090 508576 380052 508600
rect 377090 508544 379530 508576
rect 377029 508542 379530 508544
rect 97717 508539 97783 508542
rect 377029 508539 377095 508542
rect 97533 508330 97599 508333
rect 99422 508330 100004 508364
rect 97533 508328 100004 508330
rect 97533 508272 97538 508328
rect 97594 508304 100004 508328
rect 376753 508330 376819 508333
rect 379470 508330 380052 508364
rect 376753 508328 380052 508330
rect 97594 508272 99482 508304
rect 97533 508270 99482 508272
rect 376753 508272 376758 508328
rect 376814 508304 380052 508328
rect 376814 508272 379530 508304
rect 376753 508270 379530 508272
rect 97533 508267 97599 508270
rect 376753 508267 376819 508270
rect -960 501802 480 501892
rect 3325 501802 3391 501805
rect -960 501800 3391 501802
rect -960 501744 3330 501800
rect 3386 501744 3391 501800
rect -960 501742 3391 501744
rect -960 501652 480 501742
rect 3325 501739 3391 501742
rect 114318 498204 114324 498268
rect 114388 498204 114394 498268
rect 118918 498204 118924 498268
rect 118988 498204 118994 498268
rect 123334 498204 123340 498268
rect 123404 498204 123410 498268
rect 150566 498204 150572 498268
rect 150636 498204 150642 498268
rect 114326 498130 114386 498204
rect 114461 498130 114527 498133
rect 114326 498128 114527 498130
rect 114326 498072 114466 498128
rect 114522 498072 114527 498128
rect 114326 498070 114527 498072
rect 118926 498130 118986 498204
rect 123342 498133 123402 498204
rect 119337 498130 119403 498133
rect 118926 498128 119403 498130
rect 118926 498072 119342 498128
rect 119398 498072 119403 498128
rect 118926 498070 119403 498072
rect 123342 498128 123451 498133
rect 123342 498072 123390 498128
rect 123446 498072 123451 498128
rect 123342 498070 123451 498072
rect 114461 498067 114527 498070
rect 119337 498067 119403 498070
rect 123385 498067 123451 498070
rect 124806 498068 124812 498132
rect 124876 498130 124882 498132
rect 125225 498130 125291 498133
rect 124876 498128 125291 498130
rect 124876 498072 125230 498128
rect 125286 498072 125291 498128
rect 124876 498070 125291 498072
rect 124876 498068 124882 498070
rect 125225 498067 125291 498070
rect 125726 498068 125732 498132
rect 125796 498130 125802 498132
rect 126789 498130 126855 498133
rect 125796 498128 126855 498130
rect 125796 498072 126794 498128
rect 126850 498072 126855 498128
rect 125796 498070 126855 498072
rect 150574 498130 150634 498204
rect 151721 498130 151787 498133
rect 150574 498128 151787 498130
rect 150574 498072 151726 498128
rect 151782 498072 151787 498128
rect 150574 498070 151787 498072
rect 125796 498068 125802 498070
rect 126789 498067 126855 498070
rect 151721 498067 151787 498070
rect 397453 498130 397519 498133
rect 397678 498130 397684 498132
rect 397453 498128 397684 498130
rect 397453 498072 397458 498128
rect 397514 498072 397684 498128
rect 397453 498070 397684 498072
rect 397453 498067 397519 498070
rect 397678 498068 397684 498070
rect 397748 498068 397754 498132
rect 425053 498130 425119 498133
rect 425462 498130 425468 498132
rect 425053 498128 425468 498130
rect 425053 498072 425058 498128
rect 425114 498072 425468 498128
rect 425053 498070 425468 498072
rect 425053 498067 425119 498070
rect 425462 498068 425468 498070
rect 425532 498068 425538 498132
rect 583520 497844 584960 498084
rect 409873 497722 409939 497725
rect 410374 497722 410380 497724
rect 409873 497720 410380 497722
rect 409873 497664 409878 497720
rect 409934 497664 410380 497720
rect 409873 497662 410380 497664
rect 409873 497659 409939 497662
rect 410374 497660 410380 497662
rect 410444 497660 410450 497724
rect 120022 497388 120028 497452
rect 120092 497450 120098 497452
rect 121361 497450 121427 497453
rect 120092 497448 121427 497450
rect 120092 497392 121366 497448
rect 121422 497392 121427 497448
rect 120092 497390 121427 497392
rect 120092 497388 120098 497390
rect 121361 497387 121427 497390
rect 398925 497314 398991 497317
rect 399886 497314 399892 497316
rect 398925 497312 399892 497314
rect 398925 497256 398930 497312
rect 398986 497256 399892 497312
rect 398925 497254 399892 497256
rect 398925 497251 398991 497254
rect 399886 497252 399892 497254
rect 399956 497252 399962 497316
rect 403157 497314 403223 497317
rect 403382 497314 403388 497316
rect 403157 497312 403388 497314
rect 403157 497256 403162 497312
rect 403218 497256 403388 497312
rect 403157 497254 403388 497256
rect 403157 497251 403223 497254
rect 403382 497252 403388 497254
rect 403452 497252 403458 497316
rect 398833 497178 398899 497181
rect 398966 497178 398972 497180
rect 398833 497176 398972 497178
rect 398833 497120 398838 497176
rect 398894 497120 398972 497176
rect 398833 497118 398972 497120
rect 398833 497115 398899 497118
rect 398966 497116 398972 497118
rect 399036 497116 399042 497180
rect 404353 497042 404419 497045
rect 405222 497042 405228 497044
rect 404353 497040 405228 497042
rect 404353 496984 404358 497040
rect 404414 496984 405228 497040
rect 404353 496982 405228 496984
rect 404353 496979 404419 496982
rect 405222 496980 405228 496982
rect 405292 496980 405298 497044
rect 113081 496908 113147 496909
rect 115473 496908 115539 496909
rect 113030 496906 113036 496908
rect 112990 496846 113036 496906
rect 113100 496904 113147 496908
rect 115422 496906 115428 496908
rect 113142 496848 113147 496904
rect 113030 496844 113036 496846
rect 113100 496844 113147 496848
rect 115382 496846 115428 496906
rect 115492 496904 115539 496908
rect 115534 496848 115539 496904
rect 115422 496844 115428 496846
rect 115492 496844 115539 496848
rect 117630 496844 117636 496908
rect 117700 496906 117706 496908
rect 118601 496906 118667 496909
rect 117700 496904 118667 496906
rect 117700 496848 118606 496904
rect 118662 496848 118667 496904
rect 117700 496846 118667 496848
rect 117700 496844 117706 496846
rect 113081 496843 113147 496844
rect 115473 496843 115539 496844
rect 118601 496843 118667 496846
rect 121126 496844 121132 496908
rect 121196 496906 121202 496908
rect 121269 496906 121335 496909
rect 121196 496904 121335 496906
rect 121196 496848 121274 496904
rect 121330 496848 121335 496904
rect 121196 496846 121335 496848
rect 121196 496844 121202 496846
rect 121269 496843 121335 496846
rect 122414 496844 122420 496908
rect 122484 496906 122490 496908
rect 122741 496906 122807 496909
rect 122484 496904 122807 496906
rect 122484 496848 122746 496904
rect 122802 496848 122807 496904
rect 122484 496846 122807 496848
rect 122484 496844 122490 496846
rect 122741 496843 122807 496846
rect 125358 496844 125364 496908
rect 125428 496906 125434 496908
rect 125501 496906 125567 496909
rect 125428 496904 125567 496906
rect 125428 496848 125506 496904
rect 125562 496848 125567 496904
rect 125428 496846 125567 496848
rect 125428 496844 125434 496846
rect 125501 496843 125567 496846
rect 130510 496844 130516 496908
rect 130580 496906 130586 496908
rect 131021 496906 131087 496909
rect 130580 496904 131087 496906
rect 130580 496848 131026 496904
rect 131082 496848 131087 496904
rect 130580 496846 131087 496848
rect 130580 496844 130586 496846
rect 131021 496843 131087 496846
rect 135478 496844 135484 496908
rect 135548 496906 135554 496908
rect 136541 496906 136607 496909
rect 140681 496908 140747 496909
rect 140630 496906 140636 496908
rect 135548 496904 136607 496906
rect 135548 496848 136546 496904
rect 136602 496848 136607 496904
rect 135548 496846 136607 496848
rect 140590 496846 140636 496906
rect 140700 496904 140747 496908
rect 140742 496848 140747 496904
rect 135548 496844 135554 496846
rect 136541 496843 136607 496846
rect 140630 496844 140636 496846
rect 140700 496844 140747 496848
rect 145598 496844 145604 496908
rect 145668 496906 145674 496908
rect 146201 496906 146267 496909
rect 145668 496904 146267 496906
rect 145668 496848 146206 496904
rect 146262 496848 146267 496904
rect 145668 496846 146267 496848
rect 145668 496844 145674 496846
rect 140681 496843 140747 496844
rect 146201 496843 146267 496846
rect 155534 496844 155540 496908
rect 155604 496906 155610 496908
rect 155861 496906 155927 496909
rect 155604 496904 155927 496906
rect 155604 496848 155866 496904
rect 155922 496848 155927 496904
rect 155604 496846 155927 496848
rect 155604 496844 155610 496846
rect 155861 496843 155927 496846
rect 160502 496844 160508 496908
rect 160572 496906 160578 496908
rect 161381 496906 161447 496909
rect 160572 496904 161447 496906
rect 160572 496848 161386 496904
rect 161442 496848 161447 496904
rect 160572 496846 161447 496848
rect 160572 496844 160578 496846
rect 161381 496843 161447 496846
rect 391933 496906 391999 496909
rect 392894 496906 392900 496908
rect 391933 496904 392900 496906
rect 391933 496848 391938 496904
rect 391994 496848 392900 496904
rect 391933 496846 392900 496848
rect 391933 496843 391999 496846
rect 392894 496844 392900 496846
rect 392964 496844 392970 496908
rect 393313 496906 393379 496909
rect 394182 496906 394188 496908
rect 393313 496904 394188 496906
rect 393313 496848 393318 496904
rect 393374 496848 394188 496904
rect 393313 496846 394188 496848
rect 393313 496843 393379 496846
rect 394182 496844 394188 496846
rect 394252 496844 394258 496908
rect 394693 496906 394759 496909
rect 395286 496906 395292 496908
rect 394693 496904 395292 496906
rect 394693 496848 394698 496904
rect 394754 496848 395292 496904
rect 394693 496846 395292 496848
rect 394693 496843 394759 496846
rect 395286 496844 395292 496846
rect 395356 496844 395362 496908
rect 400213 496906 400279 496909
rect 400990 496906 400996 496908
rect 400213 496904 400996 496906
rect 400213 496848 400218 496904
rect 400274 496848 400996 496904
rect 400213 496846 400996 496848
rect 400213 496843 400279 496846
rect 400990 496844 400996 496846
rect 401060 496844 401066 496908
rect 401593 496906 401659 496909
rect 402094 496906 402100 496908
rect 401593 496904 402100 496906
rect 401593 496848 401598 496904
rect 401654 496848 402100 496904
rect 401593 496846 402100 496848
rect 401593 496843 401659 496846
rect 402094 496844 402100 496846
rect 402164 496844 402170 496908
rect 404445 496906 404511 496909
rect 405733 496908 405799 496909
rect 404670 496906 404676 496908
rect 404445 496904 404676 496906
rect 404445 496848 404450 496904
rect 404506 496848 404676 496904
rect 404445 496846 404676 496848
rect 404445 496843 404511 496846
rect 404670 496844 404676 496846
rect 404740 496844 404746 496908
rect 405733 496904 405780 496908
rect 405844 496906 405850 496908
rect 415393 496906 415459 496909
rect 415526 496906 415532 496908
rect 405733 496848 405738 496904
rect 405733 496844 405780 496848
rect 405844 496846 405890 496906
rect 415393 496904 415532 496906
rect 415393 496848 415398 496904
rect 415454 496848 415532 496904
rect 415393 496846 415532 496848
rect 405844 496844 405850 496846
rect 405733 496843 405799 496844
rect 415393 496843 415459 496846
rect 415526 496844 415532 496846
rect 415596 496844 415602 496908
rect 419533 496906 419599 496909
rect 420126 496906 420132 496908
rect 419533 496904 420132 496906
rect 419533 496848 419538 496904
rect 419594 496848 420132 496904
rect 419533 496846 420132 496848
rect 419533 496843 419599 496846
rect 420126 496844 420132 496846
rect 420196 496844 420202 496908
rect 429193 496906 429259 496909
rect 430430 496906 430436 496908
rect 429193 496904 430436 496906
rect 429193 496848 429198 496904
rect 429254 496848 430436 496904
rect 429193 496846 430436 496848
rect 429193 496843 429259 496846
rect 430430 496844 430436 496846
rect 430500 496844 430506 496908
rect 434713 496906 434779 496909
rect 435398 496906 435404 496908
rect 434713 496904 435404 496906
rect 434713 496848 434718 496904
rect 434774 496848 435404 496904
rect 434713 496846 435404 496848
rect 434713 496843 434779 496846
rect 435398 496844 435404 496846
rect 435468 496844 435474 496908
rect 440233 496906 440299 496909
rect 440550 496906 440556 496908
rect 440233 496904 440556 496906
rect 440233 496848 440238 496904
rect 440294 496848 440556 496904
rect 440233 496846 440556 496848
rect 440233 496843 440299 496846
rect 440550 496844 440556 496846
rect 440620 496844 440626 496908
rect -960 488596 480 488836
rect 580165 484666 580231 484669
rect 583520 484666 584960 484756
rect 580165 484664 584960 484666
rect 580165 484608 580170 484664
rect 580226 484608 584960 484664
rect 580165 484606 584960 484608
rect 580165 484603 580231 484606
rect 583520 484516 584960 484606
rect -960 475690 480 475780
rect 3325 475690 3391 475693
rect -960 475688 3391 475690
rect -960 475632 3330 475688
rect 3386 475632 3391 475688
rect -960 475630 3391 475632
rect -960 475540 480 475630
rect 3325 475627 3391 475630
rect 579981 471474 580047 471477
rect 583520 471474 584960 471564
rect 579981 471472 584960 471474
rect 579981 471416 579986 471472
rect 580042 471416 584960 471472
rect 579981 471414 584960 471416
rect 579981 471411 580047 471414
rect 583520 471324 584960 471414
rect -960 462634 480 462724
rect 3325 462634 3391 462637
rect -960 462632 3391 462634
rect -960 462576 3330 462632
rect 3386 462576 3391 462632
rect -960 462574 3391 462576
rect -960 462484 480 462574
rect 3325 462571 3391 462574
rect 580165 458146 580231 458149
rect 583520 458146 584960 458236
rect 580165 458144 584960 458146
rect 580165 458088 580170 458144
rect 580226 458088 584960 458144
rect 580165 458086 584960 458088
rect 580165 458083 580231 458086
rect 583520 457996 584960 458086
rect -960 449578 480 449668
rect 3325 449578 3391 449581
rect -960 449576 3391 449578
rect -960 449520 3330 449576
rect 3386 449520 3391 449576
rect -960 449518 3391 449520
rect -960 449428 480 449518
rect 3325 449515 3391 449518
rect 583520 444668 584960 444908
rect -960 436508 480 436748
rect 579613 431626 579679 431629
rect 583520 431626 584960 431716
rect 579613 431624 584960 431626
rect 579613 431568 579618 431624
rect 579674 431568 584960 431624
rect 579613 431566 584960 431568
rect 579613 431563 579679 431566
rect 583520 431476 584960 431566
rect -960 423602 480 423692
rect 3141 423602 3207 423605
rect -960 423600 3207 423602
rect -960 423544 3146 423600
rect 3202 423544 3207 423600
rect -960 423542 3207 423544
rect -960 423452 480 423542
rect 3141 423539 3207 423542
rect 579705 418298 579771 418301
rect 583520 418298 584960 418388
rect 579705 418296 584960 418298
rect 579705 418240 579710 418296
rect 579766 418240 584960 418296
rect 579705 418238 584960 418240
rect 579705 418235 579771 418238
rect 583520 418148 584960 418238
rect -960 410546 480 410636
rect 3141 410546 3207 410549
rect -960 410544 3207 410546
rect -960 410488 3146 410544
rect 3202 410488 3207 410544
rect -960 410486 3207 410488
rect -960 410396 480 410486
rect 3141 410483 3207 410486
rect 579981 404970 580047 404973
rect 583520 404970 584960 405060
rect 579981 404968 584960 404970
rect 579981 404912 579986 404968
rect 580042 404912 584960 404968
rect 579981 404910 584960 404912
rect 579981 404907 580047 404910
rect 583520 404820 584960 404910
rect -960 397490 480 397580
rect 3325 397490 3391 397493
rect -960 397488 3391 397490
rect -960 397432 3330 397488
rect 3386 397432 3391 397488
rect -960 397430 3391 397432
rect -960 397340 480 397430
rect 3325 397427 3391 397430
rect 4797 393954 4863 393957
rect 233785 393954 233851 393957
rect 4797 393952 233851 393954
rect 4797 393896 4802 393952
rect 4858 393896 233790 393952
rect 233846 393896 233851 393952
rect 4797 393894 233851 393896
rect 4797 393891 4863 393894
rect 233785 393891 233851 393894
rect 233785 393412 233851 393413
rect 233734 393410 233740 393412
rect 233694 393350 233740 393410
rect 233804 393408 233851 393412
rect 233846 393352 233851 393408
rect 233734 393348 233740 393350
rect 233804 393348 233851 393352
rect 233785 393347 233851 393348
rect 583520 391628 584960 391868
rect 239622 385052 239628 385116
rect 239692 385114 239698 385116
rect 270861 385114 270927 385117
rect 239692 385112 270927 385114
rect 239692 385056 270866 385112
rect 270922 385056 270927 385112
rect 239692 385054 270927 385056
rect 239692 385052 239698 385054
rect 270861 385051 270927 385054
rect 295609 384978 295675 384981
rect 295977 384978 296043 384981
rect 295609 384976 296043 384978
rect 295609 384920 295614 384976
rect 295670 384920 295982 384976
rect 296038 384920 296043 384976
rect 295609 384918 296043 384920
rect 295609 384915 295675 384918
rect 295977 384915 296043 384918
rect 273437 384842 273503 384845
rect 293350 384842 293356 384844
rect 273437 384840 293356 384842
rect 273437 384784 273442 384840
rect 273498 384784 293356 384840
rect 273437 384782 293356 384784
rect 273437 384779 273503 384782
rect 293350 384780 293356 384782
rect 293420 384780 293426 384844
rect 295333 384842 295399 384845
rect 296294 384842 296300 384844
rect 295333 384840 296300 384842
rect 295333 384784 295338 384840
rect 295394 384784 296300 384840
rect 295333 384782 296300 384784
rect 295333 384779 295399 384782
rect 296294 384780 296300 384782
rect 296364 384780 296370 384844
rect 273069 384706 273135 384709
rect 295006 384706 295012 384708
rect 273069 384704 295012 384706
rect 273069 384648 273074 384704
rect 273130 384648 295012 384704
rect 273069 384646 295012 384648
rect 273069 384643 273135 384646
rect 295006 384644 295012 384646
rect 295076 384644 295082 384708
rect -960 384284 480 384524
rect 238518 384508 238524 384572
rect 238588 384570 238594 384572
rect 281073 384570 281139 384573
rect 238588 384568 281139 384570
rect 238588 384512 281078 384568
rect 281134 384512 281139 384568
rect 238588 384510 281139 384512
rect 238588 384508 238594 384510
rect 281073 384507 281139 384510
rect 239213 384434 239279 384437
rect 267641 384434 267707 384437
rect 239213 384432 267707 384434
rect 239213 384376 239218 384432
rect 239274 384376 267646 384432
rect 267702 384376 267707 384432
rect 239213 384374 267707 384376
rect 239213 384371 239279 384374
rect 267641 384371 267707 384374
rect 268193 384434 268259 384437
rect 290774 384434 290780 384436
rect 268193 384432 290780 384434
rect 268193 384376 268198 384432
rect 268254 384376 290780 384432
rect 268193 384374 290780 384376
rect 268193 384371 268259 384374
rect 290774 384372 290780 384374
rect 290844 384372 290850 384436
rect 291837 384434 291903 384437
rect 343725 384434 343791 384437
rect 291837 384432 343791 384434
rect 291837 384376 291842 384432
rect 291898 384376 343730 384432
rect 343786 384376 343791 384432
rect 291837 384374 343791 384376
rect 291837 384371 291903 384374
rect 343725 384371 343791 384374
rect 262121 384298 262187 384301
rect 345054 384298 345060 384300
rect 262121 384296 345060 384298
rect 262121 384240 262126 384296
rect 262182 384240 345060 384296
rect 262121 384238 345060 384240
rect 262121 384235 262187 384238
rect 345054 384236 345060 384238
rect 345124 384236 345130 384300
rect 238150 384100 238156 384164
rect 238220 384162 238226 384164
rect 266445 384162 266511 384165
rect 238220 384160 266511 384162
rect 238220 384104 266450 384160
rect 266506 384104 266511 384160
rect 238220 384102 266511 384104
rect 238220 384100 238226 384102
rect 266445 384099 266511 384102
rect 290917 384162 290983 384165
rect 523677 384162 523743 384165
rect 290917 384160 523743 384162
rect 290917 384104 290922 384160
rect 290978 384104 523682 384160
rect 523738 384104 523743 384160
rect 290917 384102 523743 384104
rect 290917 384099 290983 384102
rect 523677 384099 523743 384102
rect 235206 383964 235212 384028
rect 235276 384026 235282 384028
rect 268653 384026 268719 384029
rect 235276 384024 268719 384026
rect 235276 383968 268658 384024
rect 268714 383968 268719 384024
rect 235276 383966 268719 383968
rect 235276 383964 235282 383966
rect 268653 383963 268719 383966
rect 289721 384026 289787 384029
rect 580441 384026 580507 384029
rect 289721 384024 580507 384026
rect 289721 383968 289726 384024
rect 289782 383968 580446 384024
rect 580502 383968 580507 384024
rect 289721 383966 580507 383968
rect 289721 383963 289787 383966
rect 580441 383963 580507 383966
rect 242157 383890 242223 383893
rect 580625 383890 580691 383893
rect 242157 383888 580691 383890
rect 242157 383832 242162 383888
rect 242218 383832 580630 383888
rect 580686 383832 580691 383888
rect 242157 383830 580691 383832
rect 242157 383827 242223 383830
rect 580625 383827 580691 383830
rect 287881 383754 287947 383757
rect 291326 383754 291332 383756
rect 287881 383752 291332 383754
rect 287881 383696 287886 383752
rect 287942 383696 291332 383752
rect 287881 383694 291332 383696
rect 287881 383691 287947 383694
rect 291326 383692 291332 383694
rect 291396 383692 291402 383756
rect 296621 383754 296687 383757
rect 356697 383754 356763 383757
rect 296621 383752 356763 383754
rect 296621 383696 296626 383752
rect 296682 383696 356702 383752
rect 356758 383696 356763 383752
rect 296621 383694 356763 383696
rect 296621 383691 296687 383694
rect 356697 383691 356763 383694
rect 259637 383618 259703 383621
rect 260189 383618 260255 383621
rect 259637 383616 260255 383618
rect 259637 383560 259642 383616
rect 259698 383560 260194 383616
rect 260250 383560 260255 383616
rect 259637 383558 260255 383560
rect 259637 383555 259703 383558
rect 260189 383555 260255 383558
rect 271413 383346 271479 383349
rect 296846 383346 296852 383348
rect 271413 383344 296852 383346
rect 271413 383288 271418 383344
rect 271474 383288 296852 383344
rect 271413 383286 296852 383288
rect 271413 383283 271479 383286
rect 296846 383284 296852 383286
rect 296916 383284 296922 383348
rect 243261 383210 243327 383213
rect 577865 383210 577931 383213
rect 243261 383208 577931 383210
rect 243261 383152 243266 383208
rect 243322 383152 577870 383208
rect 577926 383152 577931 383208
rect 243261 383150 577931 383152
rect 243261 383147 243327 383150
rect 577865 383147 577931 383150
rect 242433 383074 242499 383077
rect 577681 383074 577747 383077
rect 242433 383072 577747 383074
rect 242433 383016 242438 383072
rect 242494 383016 577686 383072
rect 577742 383016 577747 383072
rect 242433 383014 577747 383016
rect 242433 383011 242499 383014
rect 577681 383011 577747 383014
rect 259637 382938 259703 382941
rect 290590 382938 290596 382940
rect 259637 382936 290596 382938
rect 259637 382880 259642 382936
rect 259698 382880 290596 382936
rect 259637 382878 290596 382880
rect 259637 382875 259703 382878
rect 290590 382876 290596 382878
rect 290660 382876 290666 382940
rect 235257 382802 235323 382805
rect 267549 382802 267615 382805
rect 235257 382800 267615 382802
rect 235257 382744 235262 382800
rect 235318 382744 267554 382800
rect 267610 382744 267615 382800
rect 235257 382742 267615 382744
rect 235257 382739 235323 382742
rect 267549 382739 267615 382742
rect 291101 382802 291167 382805
rect 342294 382802 342300 382804
rect 291101 382800 342300 382802
rect 291101 382744 291106 382800
rect 291162 382744 342300 382800
rect 291101 382742 342300 382744
rect 291101 382739 291167 382742
rect 342294 382740 342300 382742
rect 342364 382740 342370 382804
rect 90357 382666 90423 382669
rect 268377 382666 268443 382669
rect 90357 382664 268443 382666
rect 90357 382608 90362 382664
rect 90418 382608 268382 382664
rect 268438 382608 268443 382664
rect 90357 382606 268443 382608
rect 90357 382603 90423 382606
rect 268377 382603 268443 382606
rect 278037 382666 278103 382669
rect 342846 382666 342852 382668
rect 278037 382664 342852 382666
rect 278037 382608 278042 382664
rect 278098 382608 342852 382664
rect 278037 382606 342852 382608
rect 278037 382603 278103 382606
rect 342846 382604 342852 382606
rect 342916 382604 342922 382668
rect 276749 382530 276815 382533
rect 293166 382530 293172 382532
rect 276749 382528 293172 382530
rect 276749 382472 276754 382528
rect 276810 382472 293172 382528
rect 276749 382470 293172 382472
rect 276749 382467 276815 382470
rect 293166 382468 293172 382470
rect 293236 382468 293242 382532
rect 241421 382394 241487 382397
rect 249057 382394 249123 382397
rect 241421 382392 249123 382394
rect 241421 382336 241426 382392
rect 241482 382336 249062 382392
rect 249118 382336 249123 382392
rect 241421 382334 249123 382336
rect 241421 382331 241487 382334
rect 249057 382331 249123 382334
rect 278405 382394 278471 382397
rect 296110 382394 296116 382396
rect 278405 382392 296116 382394
rect 278405 382336 278410 382392
rect 278466 382336 296116 382392
rect 278405 382334 296116 382336
rect 278405 382331 278471 382334
rect 296110 382332 296116 382334
rect 296180 382332 296186 382396
rect 240777 382122 240843 382125
rect 246297 382122 246363 382125
rect 240777 382120 246363 382122
rect 240777 382064 240782 382120
rect 240838 382064 246302 382120
rect 246358 382064 246363 382120
rect 240777 382062 246363 382064
rect 240777 382059 240843 382062
rect 246297 382059 246363 382062
rect 274541 382122 274607 382125
rect 283971 382124 284037 382125
rect 283966 382122 283972 382124
rect 274541 382120 282930 382122
rect 274541 382064 274546 382120
rect 274602 382064 282930 382120
rect 274541 382062 282930 382064
rect 283880 382062 283972 382122
rect 274541 382059 274607 382062
rect 239673 381986 239739 381989
rect 246021 381986 246087 381989
rect 239673 381984 246087 381986
rect 239673 381928 239678 381984
rect 239734 381928 246026 381984
rect 246082 381928 246087 381984
rect 239673 381926 246087 381928
rect 239673 381923 239739 381926
rect 246021 381923 246087 381926
rect 237230 381788 237236 381852
rect 237300 381850 237306 381852
rect 257889 381850 257955 381853
rect 237300 381848 257955 381850
rect 237300 381792 257894 381848
rect 257950 381792 257955 381848
rect 237300 381790 257955 381792
rect 237300 381788 237306 381790
rect 257889 381787 257955 381790
rect 258758 381788 258764 381852
rect 258828 381850 258834 381852
rect 269205 381850 269271 381853
rect 273897 381852 273963 381853
rect 276105 381852 276171 381853
rect 273846 381850 273852 381852
rect 258828 381848 269271 381850
rect 258828 381792 269210 381848
rect 269266 381792 269271 381848
rect 258828 381790 269271 381792
rect 273806 381790 273852 381850
rect 273916 381848 273963 381852
rect 276054 381850 276060 381852
rect 273958 381792 273963 381848
rect 258828 381788 258834 381790
rect 269205 381787 269271 381790
rect 273846 381788 273852 381790
rect 273916 381788 273963 381792
rect 276014 381790 276060 381850
rect 276124 381848 276171 381852
rect 276166 381792 276171 381848
rect 276054 381788 276060 381790
rect 276124 381788 276171 381792
rect 273897 381787 273963 381788
rect 276105 381787 276171 381788
rect 277761 381850 277827 381853
rect 282453 381852 282519 381853
rect 280286 381850 280292 381852
rect 277761 381848 280292 381850
rect 277761 381792 277766 381848
rect 277822 381792 280292 381848
rect 277761 381790 280292 381792
rect 277761 381787 277827 381790
rect 280286 381788 280292 381790
rect 280356 381788 280362 381852
rect 282453 381848 282500 381852
rect 282564 381850 282570 381852
rect 282870 381850 282930 382062
rect 283966 382060 283972 382062
rect 284036 382060 284042 382124
rect 289997 382122 290063 382125
rect 290958 382122 290964 382124
rect 289997 382120 290964 382122
rect 289997 382064 290002 382120
rect 290058 382064 290964 382120
rect 289997 382062 290964 382064
rect 283971 382059 284037 382060
rect 289997 382059 290063 382062
rect 290958 382060 290964 382062
rect 291028 382060 291034 382124
rect 293907 382122 293973 382125
rect 298134 382122 298140 382124
rect 293907 382120 298140 382122
rect 293907 382064 293912 382120
rect 293968 382064 298140 382120
rect 293907 382062 298140 382064
rect 293907 382059 293973 382062
rect 298134 382060 298140 382062
rect 298204 382060 298210 382124
rect 288525 381986 288591 381989
rect 288750 381986 288756 381988
rect 288525 381984 288756 381986
rect 288525 381928 288530 381984
rect 288586 381928 288756 381984
rect 288525 381926 288756 381928
rect 288525 381923 288591 381926
rect 288750 381924 288756 381926
rect 288820 381924 288826 381988
rect 288934 381924 288940 381988
rect 289004 381986 289010 381988
rect 289353 381986 289419 381989
rect 289004 381984 289419 381986
rect 289004 381928 289358 381984
rect 289414 381928 289419 381984
rect 289004 381926 289419 381928
rect 289004 381924 289010 381926
rect 289353 381923 289419 381926
rect 291142 381924 291148 381988
rect 291212 381986 291218 381988
rect 292113 381986 292179 381989
rect 291212 381984 292179 381986
rect 291212 381928 292118 381984
rect 292174 381928 292179 381984
rect 291212 381926 292179 381928
rect 291212 381924 291218 381926
rect 292113 381923 292179 381926
rect 293902 381924 293908 381988
rect 293972 381986 293978 381988
rect 294873 381986 294939 381989
rect 293972 381984 294939 381986
rect 293972 381928 294878 381984
rect 294934 381928 294939 381984
rect 293972 381926 294939 381928
rect 293972 381924 293978 381926
rect 294873 381923 294939 381926
rect 295701 381988 295767 381989
rect 295701 381984 295748 381988
rect 295812 381986 295818 381988
rect 296253 381986 296319 381989
rect 296478 381986 296484 381988
rect 295701 381928 295706 381984
rect 295701 381924 295748 381928
rect 295812 381926 295858 381986
rect 296253 381984 296484 381986
rect 296253 381928 296258 381984
rect 296314 381928 296484 381984
rect 296253 381926 296484 381928
rect 295812 381924 295818 381926
rect 295701 381923 295767 381924
rect 296253 381923 296319 381926
rect 296478 381924 296484 381926
rect 296548 381924 296554 381988
rect 345238 381850 345244 381852
rect 282453 381792 282458 381848
rect 282453 381788 282500 381792
rect 282564 381790 282610 381850
rect 282870 381790 345244 381850
rect 282564 381788 282570 381790
rect 345238 381788 345244 381790
rect 345308 381788 345314 381852
rect 282453 381787 282519 381788
rect 241881 381714 241947 381717
rect 347037 381714 347103 381717
rect 241881 381712 347103 381714
rect 241881 381656 241886 381712
rect 241942 381656 347042 381712
rect 347098 381656 347103 381712
rect 241881 381654 347103 381656
rect 241881 381651 241947 381654
rect 347037 381651 347103 381654
rect 246297 381578 246363 381581
rect 580206 381578 580212 381580
rect 246297 381576 580212 381578
rect 246297 381520 246302 381576
rect 246358 381520 580212 381576
rect 246297 381518 580212 381520
rect 246297 381515 246363 381518
rect 580206 381516 580212 381518
rect 580276 381516 580282 381580
rect 239949 381444 240015 381445
rect 239949 381440 239996 381444
rect 240060 381442 240066 381444
rect 240501 381442 240567 381445
rect 242382 381442 242388 381444
rect 239949 381384 239954 381440
rect 239949 381380 239996 381384
rect 240060 381382 240106 381442
rect 240501 381440 242388 381442
rect 240501 381384 240506 381440
rect 240562 381384 242388 381440
rect 240501 381382 242388 381384
rect 240060 381380 240066 381382
rect 239949 381379 240015 381380
rect 240501 381379 240567 381382
rect 242382 381380 242388 381382
rect 242452 381380 242458 381444
rect 242709 381442 242775 381445
rect 245469 381444 245535 381445
rect 242709 381440 244290 381442
rect 242709 381384 242714 381440
rect 242770 381384 244290 381440
rect 242709 381382 244290 381384
rect 242709 381379 242775 381382
rect 244230 381306 244290 381382
rect 245469 381440 245516 381444
rect 245580 381442 245586 381444
rect 246021 381442 246087 381445
rect 346894 381442 346900 381444
rect 245469 381384 245474 381440
rect 245469 381380 245516 381384
rect 245580 381382 245626 381442
rect 246021 381440 346900 381442
rect 246021 381384 246026 381440
rect 246082 381384 346900 381440
rect 246021 381382 346900 381384
rect 245580 381380 245586 381382
rect 245469 381379 245535 381380
rect 246021 381379 246087 381382
rect 346894 381380 346900 381382
rect 346964 381380 346970 381444
rect 407757 381306 407823 381309
rect 244230 381304 407823 381306
rect 244230 381248 407762 381304
rect 407818 381248 407823 381304
rect 244230 381246 407823 381248
rect 407757 381243 407823 381246
rect 3509 381170 3575 381173
rect 258758 381170 258764 381172
rect 3509 381168 258764 381170
rect 3509 381112 3514 381168
rect 3570 381112 258764 381168
rect 3509 381110 258764 381112
rect 3509 381107 3575 381110
rect 258758 381108 258764 381110
rect 258828 381108 258834 381172
rect 280286 381108 280292 381172
rect 280356 381170 280362 381172
rect 291694 381170 291700 381172
rect 280356 381110 291700 381170
rect 280356 381108 280362 381110
rect 291694 381108 291700 381110
rect 291764 381108 291770 381172
rect 242382 380972 242388 381036
rect 242452 381034 242458 381036
rect 580349 381034 580415 381037
rect 242452 381032 580415 381034
rect 242452 380976 580354 381032
rect 580410 380976 580415 381032
rect 242452 380974 580415 380976
rect 242452 380972 242458 380974
rect 580349 380971 580415 380974
rect 237046 380564 237052 380628
rect 237116 380626 237122 380628
rect 273846 380626 273852 380628
rect 237116 380566 273852 380626
rect 237116 380564 237122 380566
rect 273846 380564 273852 380566
rect 273916 380564 273922 380628
rect 283966 380564 283972 380628
rect 284036 380626 284042 380628
rect 301037 380626 301103 380629
rect 284036 380624 301103 380626
rect 284036 380568 301042 380624
rect 301098 380568 301103 380624
rect 284036 380566 301103 380568
rect 284036 380564 284042 380566
rect 301037 380563 301103 380566
rect 234337 380490 234403 380493
rect 276054 380490 276060 380492
rect 234337 380488 276060 380490
rect 234337 380432 234342 380488
rect 234398 380432 276060 380488
rect 234337 380430 276060 380432
rect 234337 380427 234403 380430
rect 276054 380428 276060 380430
rect 276124 380428 276130 380492
rect 282494 380428 282500 380492
rect 282564 380490 282570 380492
rect 301129 380490 301195 380493
rect 282564 380488 301195 380490
rect 282564 380432 301134 380488
rect 301190 380432 301195 380488
rect 282564 380430 301195 380432
rect 282564 380428 282570 380430
rect 301129 380427 301195 380430
rect 245510 380292 245516 380356
rect 245580 380354 245586 380356
rect 578141 380354 578207 380357
rect 245580 380352 578207 380354
rect 245580 380296 578146 380352
rect 578202 380296 578207 380352
rect 245580 380294 578207 380296
rect 245580 380292 245586 380294
rect 578141 380291 578207 380294
rect 239990 380156 239996 380220
rect 240060 380218 240066 380220
rect 577497 380218 577563 380221
rect 240060 380216 577563 380218
rect 240060 380160 577502 380216
rect 577558 380160 577563 380216
rect 240060 380158 577563 380160
rect 240060 380156 240066 380158
rect 577497 380155 577563 380158
rect 580165 378450 580231 378453
rect 583520 378450 584960 378540
rect 580165 378448 584960 378450
rect 580165 378392 580170 378448
rect 580226 378392 584960 378448
rect 580165 378390 584960 378392
rect 580165 378387 580231 378390
rect 583520 378300 584960 378390
rect 296110 374036 296116 374100
rect 296180 374098 296186 374100
rect 296662 374098 296668 374100
rect 296180 374038 296668 374098
rect 296180 374036 296186 374038
rect 296662 374036 296668 374038
rect 296732 374036 296738 374100
rect 296110 373900 296116 373964
rect 296180 373962 296186 373964
rect 296662 373962 296668 373964
rect 296180 373902 296668 373962
rect 296180 373900 296186 373902
rect 296662 373900 296668 373902
rect 296732 373900 296738 373964
rect -960 371378 480 371468
rect 3141 371378 3207 371381
rect -960 371376 3207 371378
rect -960 371320 3146 371376
rect 3202 371320 3207 371376
rect -960 371318 3207 371320
rect -960 371228 480 371318
rect 3141 371315 3207 371318
rect 580073 365122 580139 365125
rect 583520 365122 584960 365212
rect 580073 365120 584960 365122
rect 580073 365064 580078 365120
rect 580134 365064 584960 365120
rect 580073 365062 584960 365064
rect 580073 365059 580139 365062
rect 583520 364972 584960 365062
rect 296110 364380 296116 364444
rect 296180 364442 296186 364444
rect 296662 364442 296668 364444
rect 296180 364382 296668 364442
rect 296180 364380 296186 364382
rect 296662 364380 296668 364382
rect 296732 364380 296738 364444
rect 296110 364244 296116 364308
rect 296180 364306 296186 364308
rect 296662 364306 296668 364308
rect 296180 364246 296668 364306
rect 296180 364244 296186 364246
rect 296662 364244 296668 364246
rect 296732 364244 296738 364308
rect 238334 363428 238340 363492
rect 238404 363490 238410 363492
rect 238886 363490 238892 363492
rect 238404 363430 238892 363490
rect 238404 363428 238410 363430
rect 238886 363428 238892 363430
rect 238956 363428 238962 363492
rect -960 358458 480 358548
rect 3785 358458 3851 358461
rect -960 358456 3851 358458
rect -960 358400 3790 358456
rect 3846 358400 3851 358456
rect -960 358398 3851 358400
rect -960 358308 480 358398
rect 3785 358395 3851 358398
rect 296110 354724 296116 354788
rect 296180 354786 296186 354788
rect 296662 354786 296668 354788
rect 296180 354726 296668 354786
rect 296180 354724 296186 354726
rect 296662 354724 296668 354726
rect 296732 354724 296738 354788
rect 296110 354588 296116 354652
rect 296180 354650 296186 354652
rect 296662 354650 296668 354652
rect 296180 354590 296668 354650
rect 296180 354588 296186 354590
rect 296662 354588 296668 354590
rect 296732 354588 296738 354652
rect 579981 351930 580047 351933
rect 583520 351930 584960 352020
rect 579981 351928 584960 351930
rect 579981 351872 579986 351928
rect 580042 351872 584960 351928
rect 579981 351870 584960 351872
rect 579981 351867 580047 351870
rect 583520 351780 584960 351870
rect -960 345402 480 345492
rect 2957 345402 3023 345405
rect -960 345400 3023 345402
rect -960 345344 2962 345400
rect 3018 345344 3023 345400
rect -960 345342 3023 345344
rect -960 345252 480 345342
rect 2957 345339 3023 345342
rect 296110 345068 296116 345132
rect 296180 345130 296186 345132
rect 296662 345130 296668 345132
rect 296180 345070 296668 345130
rect 296180 345068 296186 345070
rect 296662 345068 296668 345070
rect 296732 345068 296738 345132
rect 296110 344932 296116 344996
rect 296180 344994 296186 344996
rect 296662 344994 296668 344996
rect 296180 344934 296668 344994
rect 296180 344932 296186 344934
rect 296662 344932 296668 344934
rect 296732 344932 296738 344996
rect 238886 339900 238892 339964
rect 238956 339962 238962 339964
rect 239622 339962 239628 339964
rect 238956 339902 239628 339962
rect 238956 339900 238962 339902
rect 239622 339900 239628 339902
rect 239692 339900 239698 339964
rect 583520 338452 584960 338692
rect 244641 338330 244707 338333
rect 244641 338328 246222 338330
rect 244641 338272 244646 338328
rect 244702 338272 246222 338328
rect 244641 338270 246222 338272
rect 244641 338267 244707 338270
rect 245878 338132 245884 338196
rect 245948 338194 245954 338196
rect 245948 338132 245992 338194
rect 245932 337959 245992 338132
rect 246162 337959 246222 338270
rect 254526 338194 254532 338196
rect 253982 338134 254532 338194
rect 253982 337959 254042 338134
rect 254526 338132 254532 338134
rect 254596 338132 254602 338196
rect 255630 338194 255636 338196
rect 255454 338134 255636 338194
rect 255454 337959 255514 338134
rect 255630 338132 255636 338134
rect 255700 338132 255706 338196
rect 291009 338194 291075 338197
rect 287608 338192 291075 338194
rect 287608 338136 291014 338192
rect 291070 338136 291075 338192
rect 287608 338134 291075 338136
rect 255814 338058 255820 338060
rect 255684 337998 255820 338058
rect 255684 337959 255744 337998
rect 255814 337996 255820 337998
rect 255884 337996 255890 338060
rect 266486 337996 266492 338060
rect 266556 338058 266562 338060
rect 266556 337998 266922 338058
rect 266556 337996 266562 337998
rect 245423 337956 245489 337959
rect 245791 337956 245857 337959
rect 245423 337954 245532 337956
rect 244365 337922 244431 337925
rect 245423 337922 245428 337954
rect 244365 337920 245428 337922
rect 244365 337864 244370 337920
rect 244426 337898 245428 337920
rect 245484 337898 245532 337954
rect 245748 337954 245857 337956
rect 245748 337924 245796 337954
rect 244426 337864 245532 337898
rect 244365 337862 245532 337864
rect 244365 337859 244431 337862
rect 245694 337860 245700 337924
rect 245764 337898 245796 337924
rect 245852 337898 245857 337954
rect 245764 337893 245857 337898
rect 245932 337954 246041 337959
rect 245932 337898 245980 337954
rect 246036 337898 246041 337954
rect 245932 337896 246041 337898
rect 245975 337893 246041 337896
rect 246159 337954 246225 337959
rect 246159 337898 246164 337954
rect 246220 337898 246225 337954
rect 246159 337893 246225 337898
rect 246527 337956 246593 337959
rect 246527 337954 246636 337956
rect 246527 337898 246532 337954
rect 246588 337898 246636 337954
rect 247907 337954 247973 337959
rect 246527 337893 246636 337898
rect 245764 337862 245808 337893
rect 245764 337860 245770 337862
rect 246113 337786 246179 337789
rect 246246 337786 246252 337788
rect 246113 337784 246252 337786
rect 246113 337728 246118 337784
rect 246174 337728 246252 337784
rect 246113 337726 246252 337728
rect 246113 337723 246179 337726
rect 246246 337724 246252 337726
rect 246316 337724 246322 337788
rect 244917 337650 244983 337653
rect 246576 337650 246636 337893
rect 246987 337920 247053 337925
rect 246987 337864 246992 337920
rect 247048 337864 247053 337920
rect 246987 337859 247053 337864
rect 247166 337860 247172 337924
rect 247236 337922 247242 337924
rect 247447 337922 247513 337925
rect 247236 337920 247513 337922
rect 247236 337864 247452 337920
rect 247508 337864 247513 337920
rect 247907 337898 247912 337954
rect 247968 337898 247973 337954
rect 249563 337954 249629 337959
rect 250391 337956 250457 337959
rect 247907 337893 247973 337898
rect 247236 337862 247513 337864
rect 247236 337860 247242 337862
rect 247447 337859 247513 337862
rect 246990 337789 247050 337859
rect 247910 337789 247970 337893
rect 248270 337860 248276 337924
rect 248340 337922 248346 337924
rect 248551 337922 248617 337925
rect 248340 337920 248617 337922
rect 248340 337864 248556 337920
rect 248612 337864 248617 337920
rect 249563 337898 249568 337954
rect 249624 337898 249629 337954
rect 250348 337954 250457 337956
rect 249563 337893 249629 337898
rect 249931 337922 249997 337925
rect 250110 337922 250116 337924
rect 249931 337920 250116 337922
rect 248340 337862 248617 337864
rect 248340 337860 248346 337862
rect 248551 337859 248617 337862
rect 246941 337784 247050 337789
rect 246941 337728 246946 337784
rect 247002 337728 247050 337784
rect 246941 337726 247050 337728
rect 247217 337786 247283 337789
rect 247350 337786 247356 337788
rect 247217 337784 247356 337786
rect 247217 337728 247222 337784
rect 247278 337728 247356 337784
rect 247217 337726 247356 337728
rect 246941 337723 247007 337726
rect 247217 337723 247283 337726
rect 247350 337724 247356 337726
rect 247420 337724 247426 337788
rect 247910 337784 248019 337789
rect 247910 337728 247958 337784
rect 248014 337728 248019 337784
rect 247910 337726 248019 337728
rect 247953 337723 248019 337726
rect 248689 337786 248755 337789
rect 249566 337786 249626 337893
rect 249931 337864 249936 337920
rect 249992 337864 250116 337920
rect 249931 337862 250116 337864
rect 249931 337859 249997 337862
rect 250110 337860 250116 337862
rect 250180 337860 250186 337924
rect 250348 337898 250396 337954
rect 250452 337922 250457 337954
rect 250943 337956 251009 337959
rect 250943 337954 251052 337956
rect 250452 337898 250546 337922
rect 250348 337862 250546 337898
rect 250943 337898 250948 337954
rect 251004 337898 251052 337954
rect 250943 337893 251052 337898
rect 251219 337954 251285 337959
rect 251219 337898 251224 337954
rect 251280 337922 251285 337954
rect 251955 337954 252021 337959
rect 251398 337922 251404 337924
rect 251280 337898 251404 337922
rect 251219 337893 251404 337898
rect 250207 337786 250273 337789
rect 248689 337784 249626 337786
rect 248689 337728 248694 337784
rect 248750 337728 249626 337784
rect 248689 337726 249626 337728
rect 250026 337784 250273 337786
rect 250026 337728 250212 337784
rect 250268 337728 250273 337784
rect 250026 337726 250273 337728
rect 248689 337723 248755 337726
rect 244917 337648 246636 337650
rect 244917 337592 244922 337648
rect 244978 337592 246636 337648
rect 244917 337590 246636 337592
rect 247033 337650 247099 337653
rect 249425 337650 249491 337653
rect 247033 337648 249491 337650
rect 247033 337592 247038 337648
rect 247094 337592 249430 337648
rect 249486 337592 249491 337648
rect 247033 337590 249491 337592
rect 250026 337650 250086 337726
rect 250207 337723 250273 337726
rect 250253 337650 250319 337653
rect 250486 337650 250546 337862
rect 250026 337590 250178 337650
rect 244917 337587 244983 337590
rect 247033 337587 247099 337590
rect 249425 337587 249491 337590
rect 245745 337514 245811 337517
rect 249977 337514 250043 337517
rect 245745 337512 250043 337514
rect 245745 337456 245750 337512
rect 245806 337456 249982 337512
rect 250038 337456 250043 337512
rect 245745 337454 250043 337456
rect 250118 337514 250178 337590
rect 250253 337648 250546 337650
rect 250253 337592 250258 337648
rect 250314 337592 250546 337648
rect 250253 337590 250546 337592
rect 250253 337587 250319 337590
rect 250294 337514 250300 337516
rect 250118 337454 250300 337514
rect 245745 337451 245811 337454
rect 249977 337451 250043 337454
rect 250294 337452 250300 337454
rect 250364 337452 250370 337516
rect 250805 337514 250871 337517
rect 250992 337514 251052 337893
rect 251222 337862 251404 337893
rect 251398 337860 251404 337862
rect 251468 337860 251474 337924
rect 251587 337922 251653 337925
rect 251766 337922 251772 337924
rect 251587 337920 251772 337922
rect 251587 337864 251592 337920
rect 251648 337864 251772 337920
rect 251587 337862 251772 337864
rect 251587 337859 251653 337862
rect 251766 337860 251772 337862
rect 251836 337860 251842 337924
rect 251955 337898 251960 337954
rect 252016 337898 252021 337954
rect 251955 337893 252021 337898
rect 252415 337956 252481 337959
rect 252415 337954 252616 337956
rect 252415 337898 252420 337954
rect 252476 337898 252616 337954
rect 253979 337954 254045 337959
rect 252875 337924 252941 337925
rect 252870 337922 252876 337924
rect 252415 337896 252616 337898
rect 252415 337893 252481 337896
rect 251958 337789 252018 337893
rect 251909 337784 252018 337789
rect 251909 337728 251914 337784
rect 251970 337728 252018 337784
rect 251909 337726 252018 337728
rect 252277 337786 252343 337789
rect 252556 337786 252616 337896
rect 252784 337862 252876 337922
rect 252870 337860 252876 337862
rect 252940 337860 252946 337924
rect 253059 337922 253125 337925
rect 253059 337920 253306 337922
rect 253059 337864 253064 337920
rect 253120 337864 253306 337920
rect 253979 337898 253984 337954
rect 254040 337898 254045 337954
rect 254163 337954 254229 337959
rect 254163 337924 254168 337954
rect 254224 337924 254229 337954
rect 254347 337954 254413 337959
rect 254991 337956 255057 337959
rect 253979 337893 254045 337898
rect 253059 337862 253306 337864
rect 252875 337859 252941 337860
rect 253059 337859 253125 337862
rect 253246 337789 253306 337862
rect 254158 337860 254164 337924
rect 254228 337922 254234 337924
rect 254228 337862 254286 337922
rect 254347 337898 254352 337954
rect 254408 337898 254413 337954
rect 254948 337954 255057 337956
rect 254347 337893 254413 337898
rect 254228 337860 254234 337862
rect 252783 337786 252849 337789
rect 252277 337784 252616 337786
rect 252277 337728 252282 337784
rect 252338 337728 252616 337784
rect 252277 337726 252616 337728
rect 252740 337784 252849 337786
rect 252740 337728 252788 337784
rect 252844 337728 252849 337784
rect 251909 337723 251975 337726
rect 252277 337723 252343 337726
rect 252740 337723 252849 337728
rect 253197 337784 253306 337789
rect 253197 337728 253202 337784
rect 253258 337728 253306 337784
rect 253197 337726 253306 337728
rect 253197 337723 253263 337726
rect 252740 337652 252800 337723
rect 252686 337588 252692 337652
rect 252756 337590 252800 337652
rect 252756 337588 252762 337590
rect 250805 337512 251052 337514
rect 250805 337456 250810 337512
rect 250866 337456 251052 337512
rect 250805 337454 251052 337456
rect 254350 337517 254410 337893
rect 254710 337860 254716 337924
rect 254780 337922 254786 337924
rect 254948 337922 254996 337954
rect 254780 337898 254996 337922
rect 255052 337898 255057 337954
rect 254780 337893 255057 337898
rect 255451 337954 255517 337959
rect 255451 337898 255456 337954
rect 255512 337898 255517 337954
rect 255451 337893 255517 337898
rect 255635 337954 255744 337959
rect 255635 337898 255640 337954
rect 255696 337898 255744 337954
rect 256739 337954 256805 337959
rect 255635 337896 255744 337898
rect 255819 337920 255885 337925
rect 256095 337922 256161 337925
rect 255635 337893 255701 337896
rect 254780 337862 255008 337893
rect 255819 337864 255824 337920
rect 255880 337864 255885 337920
rect 254780 337860 254786 337862
rect 255819 337859 255885 337864
rect 256052 337920 256161 337922
rect 256052 337864 256100 337920
rect 256156 337864 256161 337920
rect 256739 337898 256744 337954
rect 256800 337922 256805 337954
rect 259315 337954 259381 337959
rect 259775 337956 259841 337959
rect 257102 337922 257108 337924
rect 256800 337898 257108 337922
rect 256739 337893 257108 337898
rect 256052 337859 256161 337864
rect 256555 337886 256621 337891
rect 255543 337820 255609 337823
rect 255500 337818 255609 337820
rect 255500 337788 255548 337818
rect 255446 337724 255452 337788
rect 255516 337762 255548 337788
rect 255604 337762 255609 337818
rect 255516 337757 255609 337762
rect 255516 337726 255560 337757
rect 255516 337724 255522 337726
rect 255589 337650 255655 337653
rect 255822 337650 255882 337859
rect 255589 337648 255882 337650
rect 255589 337592 255594 337648
rect 255650 337592 255882 337648
rect 255589 337590 255882 337592
rect 255589 337587 255655 337590
rect 254350 337512 254459 337517
rect 254350 337456 254398 337512
rect 254454 337456 254459 337512
rect 254350 337454 254459 337456
rect 250805 337451 250871 337454
rect 254393 337451 254459 337454
rect 255865 337514 255931 337517
rect 256052 337514 256112 337859
rect 256555 337830 256560 337886
rect 256616 337830 256621 337886
rect 256742 337862 257108 337893
rect 257102 337860 257108 337862
rect 257172 337860 257178 337924
rect 257475 337920 257541 337925
rect 257751 337922 257817 337925
rect 257475 337864 257480 337920
rect 257536 337864 257541 337920
rect 257475 337859 257541 337864
rect 257616 337920 257817 337922
rect 257616 337864 257756 337920
rect 257812 337864 257817 337920
rect 257616 337862 257817 337864
rect 256555 337825 256621 337830
rect 256558 337653 256618 337825
rect 256509 337648 256618 337653
rect 256509 337592 256514 337648
rect 256570 337592 256618 337648
rect 256509 337590 256618 337592
rect 257478 337653 257538 337859
rect 257616 337789 257676 337862
rect 257751 337859 257817 337862
rect 258303 337922 258369 337925
rect 259126 337922 259132 337924
rect 258303 337920 259132 337922
rect 258303 337864 258308 337920
rect 258364 337864 259132 337920
rect 258303 337862 259132 337864
rect 258303 337859 258369 337862
rect 259126 337860 259132 337862
rect 259196 337860 259202 337924
rect 259315 337898 259320 337954
rect 259376 337898 259381 337954
rect 259732 337954 259841 337956
rect 259732 337924 259780 337954
rect 259315 337893 259381 337898
rect 259318 337789 259378 337893
rect 259678 337860 259684 337924
rect 259748 337898 259780 337924
rect 259836 337898 259841 337954
rect 261523 337954 261589 337959
rect 259748 337893 259841 337898
rect 260143 337922 260209 337925
rect 260971 337922 261037 337925
rect 261150 337922 261156 337924
rect 260143 337920 260482 337922
rect 259748 337862 259792 337893
rect 260143 337864 260148 337920
rect 260204 337864 260482 337920
rect 260143 337862 260482 337864
rect 259748 337860 259754 337862
rect 260143 337859 260209 337862
rect 257613 337784 257679 337789
rect 257613 337728 257618 337784
rect 257674 337728 257679 337784
rect 257613 337723 257679 337728
rect 258211 337784 258277 337789
rect 258211 337728 258216 337784
rect 258272 337728 258277 337784
rect 258211 337723 258277 337728
rect 259269 337784 259378 337789
rect 259269 337728 259274 337784
rect 259330 337728 259378 337784
rect 259269 337726 259378 337728
rect 259269 337723 259335 337726
rect 259678 337724 259684 337788
rect 259748 337786 259754 337788
rect 259867 337786 259933 337789
rect 259748 337784 259933 337786
rect 259748 337728 259872 337784
rect 259928 337728 259933 337784
rect 259748 337726 259933 337728
rect 259748 337724 259754 337726
rect 259867 337723 259933 337726
rect 257478 337648 257587 337653
rect 257478 337592 257526 337648
rect 257582 337592 257587 337648
rect 257478 337590 257587 337592
rect 256509 337587 256575 337590
rect 257521 337587 257587 337590
rect 255865 337512 256112 337514
rect 255865 337456 255870 337512
rect 255926 337456 256112 337512
rect 255865 337454 256112 337456
rect 255865 337451 255931 337454
rect 251081 337378 251147 337381
rect 251582 337378 251588 337380
rect 251081 337376 251588 337378
rect 251081 337320 251086 337376
rect 251142 337320 251588 337376
rect 251081 337318 251588 337320
rect 251081 337315 251147 337318
rect 251582 337316 251588 337318
rect 251652 337316 251658 337380
rect 253933 337378 253999 337381
rect 258214 337378 258274 337723
rect 260097 337650 260163 337653
rect 260422 337650 260482 337862
rect 260971 337920 261156 337922
rect 260971 337864 260976 337920
rect 261032 337864 261156 337920
rect 260971 337862 261156 337864
rect 260971 337859 261037 337862
rect 261150 337860 261156 337862
rect 261220 337860 261226 337924
rect 261523 337898 261528 337954
rect 261584 337898 261589 337954
rect 261523 337893 261589 337898
rect 261983 337956 262049 337959
rect 261983 337954 262092 337956
rect 261983 337898 261988 337954
rect 262044 337922 262092 337954
rect 262627 337954 262693 337959
rect 262044 337898 262184 337922
rect 261983 337893 262184 337898
rect 260097 337648 260482 337650
rect 260097 337592 260102 337648
rect 260158 337592 260482 337648
rect 260097 337590 260482 337592
rect 260097 337587 260163 337590
rect 260782 337588 260788 337652
rect 260852 337650 260858 337652
rect 261201 337650 261267 337653
rect 260852 337648 261267 337650
rect 260852 337592 261206 337648
rect 261262 337592 261267 337648
rect 260852 337590 261267 337592
rect 260852 337588 260858 337590
rect 261201 337587 261267 337590
rect 261526 337517 261586 337893
rect 262032 337862 262184 337893
rect 262124 337653 262184 337862
rect 262254 337860 262260 337924
rect 262324 337922 262330 337924
rect 262324 337860 262368 337922
rect 262438 337860 262444 337924
rect 262508 337922 262514 337924
rect 262627 337922 262632 337954
rect 262508 337898 262632 337922
rect 262688 337898 262693 337954
rect 263179 337954 263245 337959
rect 262508 337893 262693 337898
rect 262811 337920 262877 337925
rect 262508 337862 262690 337893
rect 262811 337864 262816 337920
rect 262872 337864 262877 337920
rect 263179 337898 263184 337954
rect 263240 337898 263245 337954
rect 265111 337954 265177 337959
rect 263179 337893 263245 337898
rect 263915 337922 263981 337925
rect 264094 337922 264100 337924
rect 263915 337920 264100 337922
rect 262508 337860 262514 337862
rect 262308 337789 262368 337860
rect 262811 337859 262877 337864
rect 262308 337784 262417 337789
rect 262308 337728 262356 337784
rect 262412 337728 262417 337784
rect 262308 337726 262417 337728
rect 262351 337723 262417 337726
rect 262121 337648 262187 337653
rect 262121 337592 262126 337648
rect 262182 337592 262187 337648
rect 262121 337587 262187 337592
rect 262305 337650 262371 337653
rect 262814 337650 262874 337859
rect 263041 337786 263107 337789
rect 263182 337786 263242 337893
rect 263915 337864 263920 337920
rect 263976 337864 264100 337920
rect 263915 337862 264100 337864
rect 263915 337859 263981 337862
rect 264094 337860 264100 337862
rect 264164 337860 264170 337924
rect 264467 337922 264533 337925
rect 264467 337920 264714 337922
rect 264467 337864 264472 337920
rect 264528 337864 264714 337920
rect 265111 337898 265116 337954
rect 265172 337898 265177 337954
rect 265571 337954 265637 337959
rect 265111 337893 265177 337898
rect 265387 337920 265453 337925
rect 264467 337862 264714 337864
rect 264467 337859 264533 337862
rect 264654 337789 264714 337862
rect 263731 337788 263797 337789
rect 263726 337786 263732 337788
rect 263041 337784 263242 337786
rect 263041 337728 263046 337784
rect 263102 337728 263242 337784
rect 263041 337726 263242 337728
rect 263640 337726 263732 337786
rect 263041 337723 263107 337726
rect 263726 337724 263732 337726
rect 263796 337724 263802 337788
rect 264654 337784 264763 337789
rect 264654 337728 264702 337784
rect 264758 337728 264763 337784
rect 264654 337726 264763 337728
rect 263731 337723 263797 337724
rect 264697 337723 264763 337726
rect 262305 337648 262874 337650
rect 262305 337592 262310 337648
rect 262366 337592 262874 337648
rect 262305 337590 262874 337592
rect 262305 337587 262371 337590
rect 261477 337512 261586 337517
rect 261477 337456 261482 337512
rect 261538 337456 261586 337512
rect 261477 337454 261586 337456
rect 265114 337514 265174 337893
rect 265387 337864 265392 337920
rect 265448 337864 265453 337920
rect 265571 337898 265576 337954
rect 265632 337898 265637 337954
rect 265571 337893 265637 337898
rect 266675 337920 266741 337925
rect 265387 337859 265453 337864
rect 265390 337789 265450 337859
rect 265390 337784 265499 337789
rect 265390 337728 265438 337784
rect 265494 337728 265499 337784
rect 265390 337726 265499 337728
rect 265433 337723 265499 337726
rect 265574 337653 265634 337893
rect 266123 337886 266189 337891
rect 266123 337830 266128 337886
rect 266184 337830 266189 337886
rect 266675 337864 266680 337920
rect 266736 337864 266741 337920
rect 266675 337859 266741 337864
rect 266862 337922 266922 337998
rect 270815 337954 270881 337959
rect 267595 337922 267661 337925
rect 266862 337920 267661 337922
rect 266862 337864 267600 337920
rect 267656 337864 267661 337920
rect 266862 337862 267661 337864
rect 267595 337859 267661 337862
rect 267963 337920 268029 337925
rect 267963 337864 267968 337920
rect 268024 337864 268029 337920
rect 267963 337859 268029 337864
rect 268699 337920 268765 337925
rect 268699 337864 268704 337920
rect 268760 337864 268765 337920
rect 268699 337859 268765 337864
rect 270166 337860 270172 337924
rect 270236 337922 270242 337924
rect 270447 337922 270513 337925
rect 270236 337920 270513 337922
rect 270236 337864 270452 337920
rect 270508 337864 270513 337920
rect 270815 337898 270820 337954
rect 270876 337922 270881 337954
rect 274403 337954 274469 337959
rect 272379 337924 272445 337925
rect 272374 337922 272380 337924
rect 270876 337898 272074 337922
rect 270815 337893 272074 337898
rect 270236 337862 270513 337864
rect 270818 337862 272074 337893
rect 272288 337862 272380 337922
rect 270236 337860 270242 337862
rect 270447 337859 270513 337862
rect 266123 337825 266189 337830
rect 265525 337648 265634 337653
rect 265525 337592 265530 337648
rect 265586 337592 265634 337648
rect 265525 337590 265634 337592
rect 265525 337587 265591 337590
rect 266126 337517 266186 337825
rect 266537 337650 266603 337653
rect 266678 337650 266738 337859
rect 267966 337789 268026 337859
rect 268702 337789 268762 337859
rect 267966 337784 268075 337789
rect 267966 337728 268014 337784
rect 268070 337728 268075 337784
rect 267966 337726 268075 337728
rect 268702 337784 268811 337789
rect 270401 337788 270467 337789
rect 270350 337786 270356 337788
rect 268702 337728 268750 337784
rect 268806 337728 268811 337784
rect 268702 337726 268811 337728
rect 270310 337726 270356 337786
rect 270420 337784 270467 337788
rect 271275 337786 271341 337789
rect 270462 337728 270467 337784
rect 268009 337723 268075 337726
rect 268745 337723 268811 337726
rect 270350 337724 270356 337726
rect 270420 337724 270467 337728
rect 270401 337723 270467 337724
rect 271140 337784 271341 337786
rect 271140 337728 271280 337784
rect 271336 337728 271341 337784
rect 271140 337726 271341 337728
rect 266537 337648 266738 337650
rect 266537 337592 266542 337648
rect 266598 337592 266738 337648
rect 266537 337590 266738 337592
rect 266537 337587 266603 337590
rect 271140 337517 271200 337726
rect 271275 337723 271341 337726
rect 272014 337650 272074 337862
rect 272374 337860 272380 337862
rect 272444 337860 272450 337924
rect 273667 337920 273733 337925
rect 273667 337864 273672 337920
rect 273728 337864 273733 337920
rect 272379 337859 272445 337860
rect 273667 337859 273733 337864
rect 274030 337860 274036 337924
rect 274100 337922 274106 337924
rect 274403 337922 274408 337954
rect 274100 337898 274408 337922
rect 274464 337898 274469 337954
rect 275231 337954 275297 337959
rect 274100 337893 274469 337898
rect 274587 337920 274653 337925
rect 274100 337862 274466 337893
rect 274587 337864 274592 337920
rect 274648 337864 274653 337920
rect 274100 337860 274106 337862
rect 274587 337859 274653 337864
rect 274950 337860 274956 337924
rect 275020 337922 275026 337924
rect 275231 337922 275236 337954
rect 275020 337898 275236 337922
rect 275292 337898 275297 337954
rect 277071 337954 277137 337959
rect 275020 337893 275297 337898
rect 275691 337922 275757 337925
rect 275870 337922 275876 337924
rect 275691 337920 275876 337922
rect 275020 337862 275294 337893
rect 275691 337864 275696 337920
rect 275752 337864 275876 337920
rect 275691 337862 275876 337864
rect 275020 337860 275026 337862
rect 275691 337859 275757 337862
rect 275870 337860 275876 337862
rect 275940 337860 275946 337924
rect 276054 337860 276060 337924
rect 276124 337922 276130 337924
rect 277071 337922 277076 337954
rect 276124 337898 277076 337922
rect 277132 337898 277137 337954
rect 276124 337893 277137 337898
rect 278267 337954 278333 337959
rect 278267 337898 278272 337954
rect 278328 337898 278333 337954
rect 278267 337893 278333 337898
rect 278543 337956 278609 337959
rect 278543 337954 278652 337956
rect 278543 337898 278548 337954
rect 278604 337924 278652 337954
rect 280843 337954 280909 337959
rect 278604 337898 278636 337924
rect 278543 337893 278636 337898
rect 276124 337862 277134 337893
rect 276124 337860 276130 337862
rect 272471 337786 272537 337789
rect 272471 337784 273362 337786
rect 272471 337728 272476 337784
rect 272532 337728 273362 337784
rect 272471 337726 273362 337728
rect 272471 337723 272537 337726
rect 273161 337650 273227 337653
rect 272014 337648 273227 337650
rect 272014 337592 273166 337648
rect 273222 337592 273227 337648
rect 272014 337590 273227 337592
rect 273161 337587 273227 337590
rect 265566 337514 265572 337516
rect 265114 337454 265572 337514
rect 261477 337451 261543 337454
rect 265566 337452 265572 337454
rect 265636 337452 265642 337516
rect 266077 337512 266186 337517
rect 266077 337456 266082 337512
rect 266138 337456 266186 337512
rect 266077 337454 266186 337456
rect 271137 337512 271203 337517
rect 271137 337456 271142 337512
rect 271198 337456 271203 337512
rect 266077 337451 266143 337454
rect 271137 337451 271203 337456
rect 273302 337514 273362 337726
rect 273670 337650 273730 337859
rect 274398 337724 274404 337788
rect 274468 337786 274474 337788
rect 274590 337786 274650 337859
rect 278270 337789 278330 337893
rect 278592 337862 278636 337893
rect 278630 337860 278636 337862
rect 278700 337860 278706 337924
rect 278819 337920 278885 337925
rect 278819 337864 278824 337920
rect 278880 337864 278885 337920
rect 278819 337859 278885 337864
rect 279734 337860 279740 337924
rect 279804 337922 279810 337924
rect 279923 337922 279989 337925
rect 279804 337920 279989 337922
rect 279804 337864 279928 337920
rect 279984 337864 279989 337920
rect 280383 337920 280449 337925
rect 280843 337924 280848 337954
rect 280904 337924 280909 337954
rect 286915 337954 286981 337959
rect 279804 337862 279989 337864
rect 279804 337860 279810 337862
rect 279923 337859 279989 337862
rect 280107 337886 280173 337891
rect 274468 337726 274650 337786
rect 275415 337786 275481 337789
rect 275415 337784 275938 337786
rect 275415 337728 275420 337784
rect 275476 337728 275938 337784
rect 275415 337726 275938 337728
rect 274468 337724 274474 337726
rect 275415 337723 275481 337726
rect 275878 337653 275938 337726
rect 276427 337784 276493 337789
rect 276427 337728 276432 337784
rect 276488 337728 276493 337784
rect 276427 337723 276493 337728
rect 278221 337784 278330 337789
rect 278635 337786 278701 337789
rect 278221 337728 278226 337784
rect 278282 337728 278330 337784
rect 278221 337726 278330 337728
rect 278408 337784 278701 337786
rect 278408 337728 278640 337784
rect 278696 337728 278701 337784
rect 278408 337726 278701 337728
rect 278822 337786 278882 337859
rect 280107 337830 280112 337886
rect 280168 337830 280173 337886
rect 280383 337864 280388 337920
rect 280444 337864 280449 337920
rect 280383 337859 280449 337864
rect 280838 337860 280844 337924
rect 280908 337922 280914 337924
rect 281487 337922 281553 337925
rect 282039 337922 282105 337925
rect 282315 337924 282381 337925
rect 280908 337862 280966 337922
rect 281487 337920 281688 337922
rect 281487 337864 281492 337920
rect 281548 337864 281688 337920
rect 281487 337862 281688 337864
rect 280908 337860 280914 337862
rect 281487 337859 281553 337862
rect 280107 337825 280173 337830
rect 279969 337786 280035 337789
rect 278822 337784 280035 337786
rect 278822 337728 279974 337784
rect 280030 337728 280035 337784
rect 278822 337726 280035 337728
rect 278221 337723 278287 337726
rect 273805 337650 273871 337653
rect 273670 337648 273871 337650
rect 273670 337592 273810 337648
rect 273866 337592 273871 337648
rect 273670 337590 273871 337592
rect 273805 337587 273871 337590
rect 274817 337650 274883 337653
rect 274817 337648 275018 337650
rect 274817 337592 274822 337648
rect 274878 337592 275018 337648
rect 274817 337590 275018 337592
rect 274817 337587 274883 337590
rect 274265 337514 274331 337517
rect 273302 337512 274331 337514
rect 273302 337456 274270 337512
rect 274326 337456 274331 337512
rect 273302 337454 274331 337456
rect 274265 337451 274331 337454
rect 274633 337514 274699 337517
rect 274766 337514 274772 337516
rect 274633 337512 274772 337514
rect 274633 337456 274638 337512
rect 274694 337456 274772 337512
rect 274633 337454 274772 337456
rect 274633 337451 274699 337454
rect 274766 337452 274772 337454
rect 274836 337452 274842 337516
rect 274958 337514 275018 337590
rect 275829 337648 275938 337653
rect 275829 337592 275834 337648
rect 275890 337592 275938 337648
rect 275829 337590 275938 337592
rect 276430 337653 276490 337723
rect 278408 337653 278468 337726
rect 278635 337723 278701 337726
rect 279969 337723 280035 337726
rect 276430 337648 276539 337653
rect 276430 337592 276478 337648
rect 276534 337592 276539 337648
rect 276430 337590 276539 337592
rect 275829 337587 275895 337590
rect 276473 337587 276539 337590
rect 278405 337648 278471 337653
rect 278405 337592 278410 337648
rect 278466 337592 278471 337648
rect 278405 337587 278471 337592
rect 279550 337588 279556 337652
rect 279620 337650 279626 337652
rect 280110 337650 280170 337825
rect 279620 337590 280170 337650
rect 280386 337650 280446 337859
rect 281628 337788 281688 337862
rect 282039 337920 282240 337922
rect 282039 337864 282044 337920
rect 282100 337864 282240 337920
rect 282039 337862 282240 337864
rect 282039 337859 282105 337862
rect 281574 337724 281580 337788
rect 281644 337726 281688 337788
rect 281993 337786 282059 337789
rect 282180 337786 282240 337862
rect 282310 337860 282316 337924
rect 282380 337922 282386 337924
rect 282775 337922 282841 337925
rect 283879 337922 283945 337925
rect 284431 337922 284497 337925
rect 282380 337862 282472 337922
rect 282640 337920 282841 337922
rect 282640 337864 282780 337920
rect 282836 337864 282841 337920
rect 282640 337862 282841 337864
rect 282380 337860 282386 337862
rect 282315 337859 282381 337860
rect 281993 337784 282240 337786
rect 281993 337728 281998 337784
rect 282054 337728 282240 337784
rect 281993 337726 282240 337728
rect 281644 337724 281650 337726
rect 281993 337723 282059 337726
rect 282494 337724 282500 337788
rect 282564 337786 282570 337788
rect 282640 337786 282700 337862
rect 282775 337859 282841 337862
rect 282916 337920 283945 337922
rect 282916 337864 283884 337920
rect 283940 337864 283945 337920
rect 282916 337862 283945 337864
rect 282564 337726 282700 337786
rect 282564 337724 282570 337726
rect 281349 337650 281415 337653
rect 280386 337648 281415 337650
rect 280386 337592 281354 337648
rect 281410 337592 281415 337648
rect 280386 337590 281415 337592
rect 279620 337588 279626 337590
rect 281349 337587 281415 337590
rect 282916 337517 282976 337862
rect 283879 337859 283945 337862
rect 284296 337920 284497 337922
rect 284296 337864 284436 337920
rect 284492 337864 284497 337920
rect 284296 337862 284497 337864
rect 284296 337653 284356 337862
rect 284431 337859 284497 337862
rect 284702 337860 284708 337924
rect 284772 337922 284778 337924
rect 285627 337922 285693 337925
rect 286179 337922 286245 337925
rect 284772 337920 285693 337922
rect 284772 337864 285632 337920
rect 285688 337864 285693 337920
rect 284772 337862 285693 337864
rect 284772 337860 284778 337862
rect 285627 337859 285693 337862
rect 286136 337920 286245 337922
rect 286136 337864 286184 337920
rect 286240 337864 286245 337920
rect 286136 337859 286245 337864
rect 286358 337860 286364 337924
rect 286428 337922 286434 337924
rect 286915 337922 286920 337954
rect 286428 337898 286920 337922
rect 286976 337898 286981 337954
rect 287467 337954 287533 337959
rect 286428 337893 286981 337898
rect 287283 337922 287349 337925
rect 287283 337920 287392 337922
rect 286428 337862 286978 337893
rect 287283 337864 287288 337920
rect 287344 337864 287392 337920
rect 287467 337898 287472 337954
rect 287528 337898 287533 337954
rect 287467 337893 287533 337898
rect 287608 337956 287668 338134
rect 291009 338131 291075 338134
rect 290774 337996 290780 338060
rect 290844 338058 290850 338060
rect 293953 338058 294019 338061
rect 290844 338056 294019 338058
rect 290844 338000 293958 338056
rect 294014 338000 294019 338056
rect 290844 337998 294019 338000
rect 290844 337996 290850 337998
rect 293953 337995 294019 337998
rect 287743 337956 287809 337959
rect 287608 337954 287809 337956
rect 287608 337898 287748 337954
rect 287804 337898 287809 337954
rect 287608 337896 287809 337898
rect 287743 337893 287809 337896
rect 288111 337956 288177 337959
rect 288111 337954 288220 337956
rect 288111 337898 288116 337954
rect 288172 337924 288220 337954
rect 288387 337954 288453 337959
rect 288387 337924 288392 337954
rect 288448 337924 288453 337954
rect 288939 337954 289005 337959
rect 289583 337956 289649 337959
rect 289767 337956 289833 337959
rect 290135 337956 290201 337959
rect 288172 337898 288204 337924
rect 288111 337893 288204 337898
rect 286428 337860 286434 337862
rect 287283 337859 287392 337864
rect 284983 337786 285049 337789
rect 285438 337786 285444 337788
rect 284983 337784 285444 337786
rect 284983 337728 284988 337784
rect 285044 337728 285444 337784
rect 284983 337726 285444 337728
rect 284983 337723 285049 337726
rect 285438 337724 285444 337726
rect 285508 337724 285514 337788
rect 285811 337786 285877 337789
rect 285811 337784 285920 337786
rect 285811 337728 285816 337784
rect 285872 337728 285920 337784
rect 285811 337723 285920 337728
rect 284293 337648 284359 337653
rect 284293 337592 284298 337648
rect 284354 337592 284359 337648
rect 284293 337587 284359 337592
rect 285860 337517 285920 337723
rect 286136 337517 286196 337859
rect 287332 337789 287392 337859
rect 286731 337788 286797 337789
rect 286726 337786 286732 337788
rect 286640 337726 286732 337786
rect 286726 337724 286732 337726
rect 286796 337724 286802 337788
rect 287329 337784 287395 337789
rect 287329 337728 287334 337784
rect 287390 337728 287395 337784
rect 286731 337723 286797 337724
rect 287329 337723 287395 337728
rect 287470 337653 287530 337893
rect 288160 337862 288204 337893
rect 288198 337860 288204 337862
rect 288268 337860 288274 337924
rect 288382 337860 288388 337924
rect 288452 337922 288458 337924
rect 288452 337862 288510 337922
rect 288939 337898 288944 337954
rect 289000 337898 289005 337954
rect 289540 337954 289649 337956
rect 289540 337924 289588 337954
rect 288939 337893 289005 337898
rect 288452 337860 288458 337862
rect 287830 337724 287836 337788
rect 287900 337786 287906 337788
rect 288203 337786 288269 337789
rect 287900 337784 288269 337786
rect 287900 337728 288208 337784
rect 288264 337728 288269 337784
rect 287900 337726 288269 337728
rect 287900 337724 287906 337726
rect 288203 337723 288269 337726
rect 288942 337653 289002 337893
rect 289486 337860 289492 337924
rect 289556 337898 289588 337924
rect 289644 337898 289649 337954
rect 289556 337893 289649 337898
rect 289724 337954 289833 337956
rect 289724 337898 289772 337954
rect 289828 337898 289833 337954
rect 289724 337893 289833 337898
rect 290092 337954 290201 337956
rect 290092 337898 290140 337954
rect 290196 337898 290201 337954
rect 290092 337893 290201 337898
rect 290411 337954 290477 337959
rect 290411 337898 290416 337954
rect 290472 337922 290477 337954
rect 292665 337922 292731 337925
rect 290472 337920 292731 337922
rect 290472 337898 292670 337920
rect 290411 337893 292670 337898
rect 289556 337862 289600 337893
rect 289556 337860 289562 337862
rect 289123 337784 289189 337789
rect 289123 337728 289128 337784
rect 289184 337728 289189 337784
rect 289123 337723 289189 337728
rect 289302 337724 289308 337788
rect 289372 337786 289378 337788
rect 289724 337786 289784 337893
rect 289372 337726 289784 337786
rect 290092 337786 290152 337893
rect 290414 337864 292670 337893
rect 292726 337864 292731 337920
rect 290414 337862 292731 337864
rect 292665 337859 292731 337862
rect 290273 337786 290339 337789
rect 290092 337784 290339 337786
rect 290092 337728 290278 337784
rect 290334 337728 290339 337784
rect 290092 337726 290339 337728
rect 289372 337724 289378 337726
rect 290273 337723 290339 337726
rect 287421 337648 287530 337653
rect 287421 337592 287426 337648
rect 287482 337592 287530 337648
rect 287421 337590 287530 337592
rect 288893 337648 289002 337653
rect 288893 337592 288898 337648
rect 288954 337592 289002 337648
rect 288893 337590 289002 337592
rect 287421 337587 287487 337590
rect 288893 337587 288959 337590
rect 275645 337514 275711 337517
rect 274958 337512 275711 337514
rect 274958 337456 275650 337512
rect 275706 337456 275711 337512
rect 274958 337454 275711 337456
rect 275645 337451 275711 337454
rect 282913 337512 282979 337517
rect 282913 337456 282918 337512
rect 282974 337456 282979 337512
rect 282913 337451 282979 337456
rect 285857 337512 285923 337517
rect 285857 337456 285862 337512
rect 285918 337456 285923 337512
rect 285857 337451 285923 337456
rect 286133 337512 286199 337517
rect 286133 337456 286138 337512
rect 286194 337456 286199 337512
rect 286133 337451 286199 337456
rect 288525 337514 288591 337517
rect 289126 337514 289186 337723
rect 288525 337512 289186 337514
rect 288525 337456 288530 337512
rect 288586 337456 289186 337512
rect 288525 337454 289186 337456
rect 288525 337451 288591 337454
rect 288934 337378 288940 337380
rect 253933 337376 258274 337378
rect 253933 337320 253938 337376
rect 253994 337320 258274 337376
rect 253933 337318 258274 337320
rect 273210 337318 288940 337378
rect 253933 337315 253999 337318
rect 266353 336834 266419 336837
rect 273210 336834 273270 337318
rect 288934 337316 288940 337318
rect 289004 337316 289010 337380
rect 288709 337242 288775 337245
rect 292849 337242 292915 337245
rect 288709 337240 292915 337242
rect 288709 337184 288714 337240
rect 288770 337184 292854 337240
rect 292910 337184 292915 337240
rect 288709 337182 292915 337184
rect 288709 337179 288775 337182
rect 292849 337179 292915 337182
rect 280889 336834 280955 336837
rect 266353 336832 273270 336834
rect 266353 336776 266358 336832
rect 266414 336776 273270 336832
rect 266353 336774 273270 336776
rect 280340 336832 280955 336834
rect 280340 336776 280894 336832
rect 280950 336776 280955 336832
rect 280340 336774 280955 336776
rect 266353 336771 266419 336774
rect 280340 336701 280400 336774
rect 280889 336771 280955 336774
rect 281901 336834 281967 336837
rect 283465 336836 283531 336837
rect 282678 336834 282684 336836
rect 281901 336832 282684 336834
rect 281901 336776 281906 336832
rect 281962 336776 282684 336832
rect 281901 336774 282684 336776
rect 281901 336771 281967 336774
rect 282678 336772 282684 336774
rect 282748 336772 282754 336836
rect 283414 336834 283420 336836
rect 283374 336774 283420 336834
rect 283484 336832 283531 336836
rect 283526 336776 283531 336832
rect 283414 336772 283420 336774
rect 283484 336772 283531 336776
rect 285070 336772 285076 336836
rect 285140 336834 285146 336836
rect 285305 336834 285371 336837
rect 285140 336832 285371 336834
rect 285140 336776 285310 336832
rect 285366 336776 285371 336832
rect 285140 336774 285371 336776
rect 285140 336772 285146 336774
rect 283465 336771 283531 336772
rect 285305 336771 285371 336774
rect 245561 336698 245627 336701
rect 253197 336698 253263 336701
rect 245561 336696 253263 336698
rect 245561 336640 245566 336696
rect 245622 336640 253202 336696
rect 253258 336640 253263 336696
rect 245561 336638 253263 336640
rect 245561 336635 245627 336638
rect 253197 336635 253263 336638
rect 263869 336700 263935 336701
rect 263869 336696 263916 336700
rect 263980 336698 263986 336700
rect 263869 336640 263874 336696
rect 263869 336636 263916 336640
rect 263980 336638 264026 336698
rect 263980 336636 263986 336638
rect 266302 336636 266308 336700
rect 266372 336698 266378 336700
rect 267457 336698 267523 336701
rect 266372 336696 267523 336698
rect 266372 336640 267462 336696
rect 267518 336640 267523 336696
rect 266372 336638 267523 336640
rect 266372 336636 266378 336638
rect 263869 336635 263935 336636
rect 267457 336635 267523 336638
rect 280337 336696 280403 336701
rect 280889 336700 280955 336701
rect 280337 336640 280342 336696
rect 280398 336640 280403 336696
rect 280337 336635 280403 336640
rect 280838 336636 280844 336700
rect 280908 336698 280955 336700
rect 283189 336698 283255 336701
rect 290089 336698 290155 336701
rect 280908 336696 281000 336698
rect 280950 336640 281000 336696
rect 280908 336638 281000 336640
rect 283189 336696 290155 336698
rect 283189 336640 283194 336696
rect 283250 336640 290094 336696
rect 290150 336640 290155 336696
rect 283189 336638 290155 336640
rect 280908 336636 280955 336638
rect 280889 336635 280955 336636
rect 283189 336635 283255 336638
rect 290089 336635 290155 336638
rect 292665 336698 292731 336701
rect 311157 336698 311223 336701
rect 292665 336696 311223 336698
rect 292665 336640 292670 336696
rect 292726 336640 311162 336696
rect 311218 336640 311223 336696
rect 292665 336638 311223 336640
rect 292665 336635 292731 336638
rect 311157 336635 311223 336638
rect 258022 336500 258028 336564
rect 258092 336562 258098 336564
rect 258349 336562 258415 336565
rect 258092 336560 258415 336562
rect 258092 336504 258354 336560
rect 258410 336504 258415 336560
rect 258092 336502 258415 336504
rect 258092 336500 258098 336502
rect 258349 336499 258415 336502
rect 281574 336500 281580 336564
rect 281644 336562 281650 336564
rect 382917 336562 382983 336565
rect 281644 336560 382983 336562
rect 281644 336504 382922 336560
rect 382978 336504 382983 336560
rect 281644 336502 382983 336504
rect 281644 336500 281650 336502
rect 382917 336499 382983 336502
rect 182817 336426 182883 336429
rect 245009 336426 245075 336429
rect 182817 336424 245075 336426
rect 182817 336368 182822 336424
rect 182878 336368 245014 336424
rect 245070 336368 245075 336424
rect 182817 336366 245075 336368
rect 182817 336363 182883 336366
rect 245009 336363 245075 336366
rect 285438 336364 285444 336428
rect 285508 336426 285514 336428
rect 285581 336426 285647 336429
rect 285508 336424 285647 336426
rect 285508 336368 285586 336424
rect 285642 336368 285647 336424
rect 285508 336366 285647 336368
rect 285508 336364 285514 336366
rect 285581 336363 285647 336366
rect 287605 336426 287671 336429
rect 474733 336426 474799 336429
rect 287605 336424 474799 336426
rect 287605 336368 287610 336424
rect 287666 336368 474738 336424
rect 474794 336368 474799 336424
rect 287605 336366 474799 336368
rect 287605 336363 287671 336366
rect 474733 336363 474799 336366
rect 178861 336290 178927 336293
rect 245101 336290 245167 336293
rect 254158 336290 254164 336292
rect 178861 336288 245167 336290
rect 178861 336232 178866 336288
rect 178922 336232 245106 336288
rect 245162 336232 245167 336288
rect 178861 336230 245167 336232
rect 178861 336227 178927 336230
rect 245101 336227 245167 336230
rect 245886 336230 254164 336290
rect 178677 336154 178743 336157
rect 244641 336154 244707 336157
rect 178677 336152 244707 336154
rect 178677 336096 178682 336152
rect 178738 336096 244646 336152
rect 244702 336096 244707 336152
rect 178677 336094 244707 336096
rect 178677 336091 178743 336094
rect 244641 336091 244707 336094
rect 245469 336154 245535 336157
rect 245886 336154 245946 336230
rect 254158 336228 254164 336230
rect 254228 336228 254234 336292
rect 262622 336228 262628 336292
rect 262692 336290 262698 336292
rect 271689 336290 271755 336293
rect 262692 336288 271755 336290
rect 262692 336232 271694 336288
rect 271750 336232 271755 336288
rect 262692 336230 271755 336232
rect 262692 336228 262698 336230
rect 271689 336227 271755 336230
rect 279877 336290 279943 336293
rect 280705 336290 280771 336293
rect 279877 336288 280771 336290
rect 279877 336232 279882 336288
rect 279938 336232 280710 336288
rect 280766 336232 280771 336288
rect 279877 336230 280771 336232
rect 279877 336227 279943 336230
rect 280705 336227 280771 336230
rect 282729 336290 282795 336293
rect 480253 336290 480319 336293
rect 282729 336288 480319 336290
rect 282729 336232 282734 336288
rect 282790 336232 480258 336288
rect 480314 336232 480319 336288
rect 282729 336230 480319 336232
rect 282729 336227 282795 336230
rect 480253 336227 480319 336230
rect 245469 336152 245946 336154
rect 245469 336096 245474 336152
rect 245530 336096 245946 336152
rect 245469 336094 245946 336096
rect 246849 336154 246915 336157
rect 258257 336154 258323 336157
rect 272425 336156 272491 336157
rect 246849 336152 258323 336154
rect 246849 336096 246854 336152
rect 246910 336096 258262 336152
rect 258318 336096 258323 336152
rect 246849 336094 258323 336096
rect 245469 336091 245535 336094
rect 246849 336091 246915 336094
rect 258257 336091 258323 336094
rect 272374 336092 272380 336156
rect 272444 336154 272491 336156
rect 285765 336154 285831 336157
rect 290089 336154 290155 336157
rect 487153 336154 487219 336157
rect 272444 336152 272536 336154
rect 272486 336096 272536 336152
rect 272444 336094 272536 336096
rect 285765 336152 289186 336154
rect 285765 336096 285770 336152
rect 285826 336096 289186 336152
rect 285765 336094 289186 336096
rect 272444 336092 272491 336094
rect 272425 336091 272491 336092
rect 285765 336091 285831 336094
rect 164233 336018 164299 336021
rect 258073 336018 258139 336021
rect 164233 336016 258139 336018
rect 164233 335960 164238 336016
rect 164294 335960 258078 336016
rect 258134 335960 258139 336016
rect 164233 335958 258139 335960
rect 164233 335955 164299 335958
rect 258073 335955 258139 335958
rect 277117 336020 277183 336021
rect 277117 336016 277164 336020
rect 277228 336018 277234 336020
rect 277117 335960 277122 336016
rect 277117 335956 277164 335960
rect 277228 335958 277274 336018
rect 277228 335956 277234 335958
rect 282310 335956 282316 336020
rect 282380 336018 282386 336020
rect 287605 336018 287671 336021
rect 282380 336016 287671 336018
rect 282380 335960 287610 336016
rect 287666 335960 287671 336016
rect 282380 335958 287671 335960
rect 289126 336018 289186 336094
rect 290089 336152 487219 336154
rect 290089 336096 290094 336152
rect 290150 336096 487158 336152
rect 487214 336096 487219 336152
rect 290089 336094 487219 336096
rect 290089 336091 290155 336094
rect 487153 336091 487219 336094
rect 518893 336018 518959 336021
rect 289126 336016 518959 336018
rect 289126 335960 518898 336016
rect 518954 335960 518959 336016
rect 289126 335958 518959 335960
rect 282380 335956 282386 335958
rect 277117 335955 277183 335956
rect 287605 335955 287671 335958
rect 518893 335955 518959 335958
rect 245009 335882 245075 335885
rect 254710 335882 254716 335884
rect 245009 335880 254716 335882
rect 245009 335824 245014 335880
rect 245070 335824 254716 335880
rect 245009 335822 254716 335824
rect 245009 335819 245075 335822
rect 254710 335820 254716 335822
rect 254780 335820 254786 335884
rect 255262 335820 255268 335884
rect 255332 335882 255338 335884
rect 255957 335882 256023 335885
rect 255332 335880 256023 335882
rect 255332 335824 255962 335880
rect 256018 335824 256023 335880
rect 255332 335822 256023 335824
rect 255332 335820 255338 335822
rect 255957 335819 256023 335822
rect 258165 335882 258231 335885
rect 259494 335882 259500 335884
rect 258165 335880 259500 335882
rect 258165 335824 258170 335880
rect 258226 335824 259500 335880
rect 258165 335822 259500 335824
rect 258165 335819 258231 335822
rect 259494 335820 259500 335822
rect 259564 335820 259570 335884
rect 262438 335820 262444 335884
rect 262508 335882 262514 335884
rect 262581 335882 262647 335885
rect 262508 335880 262647 335882
rect 262508 335824 262586 335880
rect 262642 335824 262647 335880
rect 262508 335822 262647 335824
rect 262508 335820 262514 335822
rect 262581 335819 262647 335822
rect 283598 335820 283604 335884
rect 283668 335882 283674 335884
rect 284017 335882 284083 335885
rect 283668 335880 284083 335882
rect 283668 335824 284022 335880
rect 284078 335824 284083 335880
rect 283668 335822 284083 335824
rect 283668 335820 283674 335822
rect 284017 335819 284083 335822
rect 243813 335746 243879 335749
rect 245561 335746 245627 335749
rect 243813 335744 245627 335746
rect 243813 335688 243818 335744
rect 243874 335688 245566 335744
rect 245622 335688 245627 335744
rect 243813 335686 245627 335688
rect 243813 335683 243879 335686
rect 245561 335683 245627 335686
rect 259545 335746 259611 335749
rect 259862 335746 259868 335748
rect 259545 335744 259868 335746
rect 259545 335688 259550 335744
rect 259606 335688 259868 335744
rect 259545 335686 259868 335688
rect 259545 335683 259611 335686
rect 259862 335684 259868 335686
rect 259932 335684 259938 335748
rect 268142 335684 268148 335748
rect 268212 335746 268218 335748
rect 269021 335746 269087 335749
rect 268212 335744 269087 335746
rect 268212 335688 269026 335744
rect 269082 335688 269087 335744
rect 268212 335686 269087 335688
rect 268212 335684 268218 335686
rect 269021 335683 269087 335686
rect 280981 335746 281047 335749
rect 280981 335744 292590 335746
rect 280981 335688 280986 335744
rect 281042 335688 292590 335744
rect 280981 335686 292590 335688
rect 280981 335683 281047 335686
rect 245377 335610 245443 335613
rect 265249 335612 265315 335613
rect 248270 335610 248276 335612
rect 245377 335608 248276 335610
rect 245377 335552 245382 335608
rect 245438 335552 248276 335608
rect 245377 335550 248276 335552
rect 245377 335547 245443 335550
rect 248270 335548 248276 335550
rect 248340 335548 248346 335612
rect 265198 335610 265204 335612
rect 265158 335550 265204 335610
rect 265268 335608 265315 335612
rect 265310 335552 265315 335608
rect 265198 335548 265204 335550
rect 265268 335548 265315 335552
rect 268326 335548 268332 335612
rect 268396 335610 268402 335612
rect 268837 335610 268903 335613
rect 268396 335608 268903 335610
rect 268396 335552 268842 335608
rect 268898 335552 268903 335608
rect 268396 335550 268903 335552
rect 268396 335548 268402 335550
rect 265249 335547 265315 335548
rect 268837 335547 268903 335550
rect 283782 335548 283788 335612
rect 283852 335610 283858 335612
rect 284201 335610 284267 335613
rect 283852 335608 284267 335610
rect 283852 335552 284206 335608
rect 284262 335552 284267 335608
rect 283852 335550 284267 335552
rect 283852 335548 283858 335550
rect 284201 335547 284267 335550
rect 284886 335548 284892 335612
rect 284956 335610 284962 335612
rect 285489 335610 285555 335613
rect 284956 335608 285555 335610
rect 284956 335552 285494 335608
rect 285550 335552 285555 335608
rect 284956 335550 285555 335552
rect 284956 335548 284962 335550
rect 285489 335547 285555 335550
rect 242525 335474 242591 335477
rect 245469 335474 245535 335477
rect 265065 335476 265131 335477
rect 265433 335476 265499 335477
rect 265014 335474 265020 335476
rect 242525 335472 245535 335474
rect 242525 335416 242530 335472
rect 242586 335416 245474 335472
rect 245530 335416 245535 335472
rect 242525 335414 245535 335416
rect 264974 335414 265020 335474
rect 265084 335472 265131 335476
rect 265382 335474 265388 335476
rect 265126 335416 265131 335472
rect 242525 335411 242591 335414
rect 245469 335411 245535 335414
rect 265014 335412 265020 335414
rect 265084 335412 265131 335416
rect 265342 335414 265388 335474
rect 265452 335472 265499 335476
rect 265494 335416 265499 335472
rect 265382 335412 265388 335414
rect 265452 335412 265499 335416
rect 268510 335412 268516 335476
rect 268580 335474 268586 335476
rect 268929 335474 268995 335477
rect 268580 335472 268995 335474
rect 268580 335416 268934 335472
rect 268990 335416 268995 335472
rect 268580 335414 268995 335416
rect 268580 335412 268586 335414
rect 265065 335411 265131 335412
rect 265433 335411 265499 335412
rect 268929 335411 268995 335414
rect 269062 335412 269068 335476
rect 269132 335474 269138 335476
rect 269481 335474 269547 335477
rect 269132 335472 269547 335474
rect 269132 335416 269486 335472
rect 269542 335416 269547 335472
rect 269132 335414 269547 335416
rect 269132 335412 269138 335414
rect 269481 335411 269547 335414
rect 271638 335412 271644 335476
rect 271708 335474 271714 335476
rect 271781 335474 271847 335477
rect 283465 335476 283531 335477
rect 283414 335474 283420 335476
rect 271708 335472 271847 335474
rect 271708 335416 271786 335472
rect 271842 335416 271847 335472
rect 271708 335414 271847 335416
rect 283374 335414 283420 335474
rect 283484 335472 283531 335476
rect 283925 335476 283991 335477
rect 284109 335476 284175 335477
rect 283925 335474 283972 335476
rect 283526 335416 283531 335472
rect 271708 335412 271714 335414
rect 271781 335411 271847 335414
rect 283414 335412 283420 335414
rect 283484 335412 283531 335416
rect 283880 335472 283972 335474
rect 283880 335416 283930 335472
rect 283880 335414 283972 335416
rect 283465 335411 283531 335412
rect 283925 335412 283972 335414
rect 284036 335412 284042 335476
rect 284109 335472 284156 335476
rect 284220 335474 284226 335476
rect 285305 335474 285371 335477
rect 290641 335474 290707 335477
rect 284109 335416 284114 335472
rect 284109 335412 284156 335416
rect 284220 335414 284266 335474
rect 285305 335472 286610 335474
rect 285305 335416 285310 335472
rect 285366 335416 286610 335472
rect 285305 335414 286610 335416
rect 284220 335412 284226 335414
rect 283925 335411 283991 335412
rect 284109 335411 284175 335412
rect 285305 335411 285371 335414
rect 243486 335276 243492 335340
rect 243556 335338 243562 335340
rect 247125 335338 247191 335341
rect 243556 335336 247191 335338
rect 243556 335280 247130 335336
rect 247186 335280 247191 335336
rect 243556 335278 247191 335280
rect 243556 335276 243562 335278
rect 247125 335275 247191 335278
rect 256918 335276 256924 335340
rect 256988 335338 256994 335340
rect 257061 335338 257127 335341
rect 261017 335340 261083 335341
rect 260966 335338 260972 335340
rect 256988 335336 257127 335338
rect 256988 335280 257066 335336
rect 257122 335280 257127 335336
rect 256988 335278 257127 335280
rect 260926 335278 260972 335338
rect 261036 335336 261083 335340
rect 261078 335280 261083 335336
rect 256988 335276 256994 335278
rect 257061 335275 257127 335278
rect 260966 335276 260972 335278
rect 261036 335276 261083 335280
rect 261017 335275 261083 335276
rect 274633 335338 274699 335341
rect 275001 335340 275067 335341
rect 274766 335338 274772 335340
rect 274633 335336 274772 335338
rect 274633 335280 274638 335336
rect 274694 335280 274772 335336
rect 274633 335278 274772 335280
rect 274633 335275 274699 335278
rect 274766 335276 274772 335278
rect 274836 335276 274842 335340
rect 274950 335276 274956 335340
rect 275020 335338 275067 335340
rect 286550 335338 286610 335414
rect 286918 335414 287898 335474
rect 286918 335338 286978 335414
rect 275020 335336 275112 335338
rect 275062 335280 275112 335336
rect 275020 335278 275112 335280
rect 286550 335278 286978 335338
rect 287838 335338 287898 335414
rect 289862 335472 290707 335474
rect 289862 335416 290646 335472
rect 290702 335416 290707 335472
rect 289862 335414 290707 335416
rect 292530 335474 292590 335686
rect 295977 335474 296043 335477
rect 292530 335472 296043 335474
rect 292530 335416 295982 335472
rect 296038 335416 296043 335472
rect 292530 335414 296043 335416
rect 289862 335338 289922 335414
rect 290641 335411 290707 335414
rect 295977 335411 296043 335414
rect 296110 335412 296116 335476
rect 296180 335474 296186 335476
rect 296662 335474 296668 335476
rect 296180 335414 296668 335474
rect 296180 335412 296186 335414
rect 296662 335412 296668 335414
rect 296732 335412 296738 335476
rect 296621 335338 296687 335341
rect 287838 335278 289922 335338
rect 296576 335336 296730 335338
rect 296576 335280 296626 335336
rect 296682 335280 296730 335336
rect 296576 335278 296730 335280
rect 275020 335276 275067 335278
rect 275001 335275 275067 335276
rect 296621 335275 296730 335278
rect 286869 335204 286935 335205
rect 296670 335204 296730 335275
rect 286869 335200 286916 335204
rect 286980 335202 286986 335204
rect 286869 335144 286874 335200
rect 286869 335140 286916 335144
rect 286980 335142 287026 335202
rect 286980 335140 286986 335142
rect 296662 335140 296668 335204
rect 296732 335140 296738 335204
rect 286869 335139 286935 335140
rect 289302 335004 289308 335068
rect 289372 335066 289378 335068
rect 289721 335066 289787 335069
rect 289372 335064 289787 335066
rect 289372 335008 289726 335064
rect 289782 335008 289787 335064
rect 289372 335006 289787 335008
rect 289372 335004 289378 335006
rect 289721 335003 289787 335006
rect 245929 334794 245995 334797
rect 246062 334794 246068 334796
rect 245929 334792 246068 334794
rect 245929 334736 245934 334792
rect 245990 334736 246068 334792
rect 245929 334734 246068 334736
rect 245929 334731 245995 334734
rect 246062 334732 246068 334734
rect 246132 334732 246138 334796
rect 252502 334732 252508 334796
rect 252572 334794 252578 334796
rect 252645 334794 252711 334797
rect 252572 334792 252711 334794
rect 252572 334736 252650 334792
rect 252706 334736 252711 334792
rect 252572 334734 252711 334736
rect 252572 334732 252578 334734
rect 252645 334731 252711 334734
rect 256734 334732 256740 334796
rect 256804 334794 256810 334796
rect 257337 334794 257403 334797
rect 256804 334792 257403 334794
rect 256804 334736 257342 334792
rect 257398 334736 257403 334792
rect 256804 334734 257403 334736
rect 256804 334732 256810 334734
rect 257337 334731 257403 334734
rect 285213 334794 285279 334797
rect 516133 334794 516199 334797
rect 285213 334792 516199 334794
rect 285213 334736 285218 334792
rect 285274 334736 516138 334792
rect 516194 334736 516199 334792
rect 285213 334734 516199 334736
rect 285213 334731 285279 334734
rect 516133 334731 516199 334734
rect 147673 334658 147739 334661
rect 256785 334658 256851 334661
rect 147673 334656 256851 334658
rect 147673 334600 147678 334656
rect 147734 334600 256790 334656
rect 256846 334600 256851 334656
rect 147673 334598 256851 334600
rect 147673 334595 147739 334598
rect 256785 334595 256851 334598
rect 288249 334658 288315 334661
rect 552013 334658 552079 334661
rect 288249 334656 552079 334658
rect 288249 334600 288254 334656
rect 288310 334600 552018 334656
rect 552074 334600 552079 334656
rect 288249 334598 552079 334600
rect 288249 334595 288315 334598
rect 552013 334595 552079 334598
rect 254117 334522 254183 334525
rect 254894 334522 254900 334524
rect 254117 334520 254900 334522
rect 254117 334464 254122 334520
rect 254178 334464 254900 334520
rect 254117 334462 254900 334464
rect 254117 334459 254183 334462
rect 254894 334460 254900 334462
rect 254964 334460 254970 334524
rect 259494 334460 259500 334524
rect 259564 334522 259570 334524
rect 259637 334522 259703 334525
rect 259564 334520 259703 334522
rect 259564 334464 259642 334520
rect 259698 334464 259703 334520
rect 259564 334462 259703 334464
rect 259564 334460 259570 334462
rect 259637 334459 259703 334462
rect 257613 333978 257679 333981
rect 291326 333978 291332 333980
rect 257613 333976 291332 333978
rect 257613 333920 257618 333976
rect 257674 333920 291332 333976
rect 257613 333918 291332 333920
rect 257613 333915 257679 333918
rect 291326 333916 291332 333918
rect 291396 333916 291402 333980
rect 282453 333842 282519 333845
rect 344502 333842 344508 333844
rect 282453 333840 344508 333842
rect 282453 333784 282458 333840
rect 282514 333784 344508 333840
rect 282453 333782 344508 333784
rect 282453 333779 282519 333782
rect 344502 333780 344508 333782
rect 344572 333780 344578 333844
rect 276565 333706 276631 333709
rect 391933 333706 391999 333709
rect 276565 333704 391999 333706
rect 276565 333648 276570 333704
rect 276626 333648 391938 333704
rect 391994 333648 391999 333704
rect 276565 333646 391999 333648
rect 276565 333643 276631 333646
rect 391933 333643 391999 333646
rect 278405 333570 278471 333573
rect 427813 333570 427879 333573
rect 278405 333568 427879 333570
rect 278405 333512 278410 333568
rect 278466 333512 427818 333568
rect 427874 333512 427879 333568
rect 278405 333510 427879 333512
rect 278405 333507 278471 333510
rect 427813 333507 427879 333510
rect 93853 333434 93919 333437
rect 251449 333434 251515 333437
rect 93853 333432 251515 333434
rect 93853 333376 93858 333432
rect 93914 333376 251454 333432
rect 251510 333376 251515 333432
rect 93853 333374 251515 333376
rect 93853 333371 93919 333374
rect 251449 333371 251515 333374
rect 279785 333434 279851 333437
rect 445753 333434 445819 333437
rect 279785 333432 445819 333434
rect 279785 333376 279790 333432
rect 279846 333376 445758 333432
rect 445814 333376 445819 333432
rect 279785 333374 445819 333376
rect 279785 333371 279851 333374
rect 445753 333371 445819 333374
rect 24853 333298 24919 333301
rect 247309 333298 247375 333301
rect 24853 333296 247375 333298
rect 24853 333240 24858 333296
rect 24914 333240 247314 333296
rect 247370 333240 247375 333296
rect 24853 333238 247375 333240
rect 24853 333235 24919 333238
rect 247309 333235 247375 333238
rect 248505 333298 248571 333301
rect 251265 333300 251331 333301
rect 248638 333298 248644 333300
rect 248505 333296 248644 333298
rect 248505 333240 248510 333296
rect 248566 333240 248644 333296
rect 248505 333238 248644 333240
rect 248505 333235 248571 333238
rect 248638 333236 248644 333238
rect 248708 333236 248714 333300
rect 251214 333236 251220 333300
rect 251284 333298 251331 333300
rect 251284 333296 251376 333298
rect 251326 333240 251376 333296
rect 251284 333238 251376 333240
rect 251284 333236 251331 333238
rect 274214 333236 274220 333300
rect 274284 333298 274290 333300
rect 274449 333298 274515 333301
rect 278497 333300 278563 333301
rect 274284 333296 274515 333298
rect 274284 333240 274454 333296
rect 274510 333240 274515 333296
rect 274284 333238 274515 333240
rect 274284 333236 274290 333238
rect 251265 333235 251331 333236
rect 274449 333235 274515 333238
rect 278446 333236 278452 333300
rect 278516 333298 278563 333300
rect 280797 333298 280863 333301
rect 463693 333298 463759 333301
rect 278516 333296 278608 333298
rect 278558 333240 278608 333296
rect 278516 333238 278608 333240
rect 280797 333296 463759 333298
rect 280797 333240 280802 333296
rect 280858 333240 463698 333296
rect 463754 333240 463759 333296
rect 280797 333238 463759 333240
rect 278516 333236 278563 333238
rect 278497 333235 278563 333236
rect 280797 333235 280863 333238
rect 463693 333235 463759 333238
rect 247401 333162 247467 333165
rect 248822 333162 248828 333164
rect 247401 333160 248828 333162
rect 247401 333104 247406 333160
rect 247462 333104 248828 333160
rect 247401 333102 248828 333104
rect 247401 333099 247467 333102
rect 248822 333100 248828 333102
rect 248892 333100 248898 333164
rect 254209 332890 254275 332893
rect 254710 332890 254716 332892
rect 254209 332888 254716 332890
rect 254209 332832 254214 332888
rect 254270 332832 254716 332888
rect 254209 332830 254716 332832
rect 254209 332827 254275 332830
rect 254710 332828 254716 332830
rect 254780 332828 254786 332892
rect -960 332196 480 332436
rect 257889 332210 257955 332213
rect 298134 332210 298140 332212
rect 257889 332208 298140 332210
rect 257889 332152 257894 332208
rect 257950 332152 298140 332208
rect 257889 332150 298140 332152
rect 257889 332147 257955 332150
rect 298134 332148 298140 332150
rect 298204 332148 298210 332212
rect 291193 332074 291259 332077
rect 535453 332074 535519 332077
rect 291193 332072 535519 332074
rect 291193 332016 291198 332072
rect 291254 332016 535458 332072
rect 535514 332016 535519 332072
rect 291193 332014 535519 332016
rect 291193 332011 291259 332014
rect 535453 332011 535519 332014
rect 243537 331938 243603 331941
rect 260782 331938 260788 331940
rect 243537 331936 260788 331938
rect 243537 331880 243542 331936
rect 243598 331880 260788 331936
rect 243537 331878 260788 331880
rect 243537 331875 243603 331878
rect 260782 331876 260788 331878
rect 260852 331876 260858 331940
rect 288198 331876 288204 331940
rect 288268 331938 288274 331940
rect 549253 331938 549319 331941
rect 288268 331936 549319 331938
rect 288268 331880 549258 331936
rect 549314 331880 549319 331936
rect 288268 331878 549319 331880
rect 288268 331876 288274 331878
rect 549253 331875 549319 331878
rect 45553 331802 45619 331805
rect 248965 331802 249031 331805
rect 45553 331800 249031 331802
rect 45553 331744 45558 331800
rect 45614 331744 248970 331800
rect 249026 331744 249031 331800
rect 45553 331742 249031 331744
rect 45553 331739 45619 331742
rect 248965 331739 249031 331742
rect 289118 331740 289124 331804
rect 289188 331802 289194 331804
rect 571333 331802 571399 331805
rect 289188 331800 571399 331802
rect 289188 331744 571338 331800
rect 571394 331744 571399 331800
rect 289188 331742 571399 331744
rect 289188 331740 289194 331742
rect 571333 331739 571399 331742
rect 263542 331196 263548 331260
rect 263612 331258 263618 331260
rect 264094 331258 264100 331260
rect 263612 331198 264100 331258
rect 263612 331196 263618 331198
rect 264094 331196 264100 331198
rect 264164 331196 264170 331260
rect 263501 331124 263567 331125
rect 263501 331122 263548 331124
rect 263456 331120 263548 331122
rect 263456 331064 263506 331120
rect 263456 331062 263548 331064
rect 263501 331060 263548 331062
rect 263612 331060 263618 331124
rect 263501 331059 263567 331060
rect 146293 330578 146359 330581
rect 257102 330578 257108 330580
rect 146293 330576 257108 330578
rect 146293 330520 146298 330576
rect 146354 330520 257108 330576
rect 146293 330518 257108 330520
rect 146293 330515 146359 330518
rect 257102 330516 257108 330518
rect 257172 330516 257178 330580
rect 284150 330516 284156 330580
rect 284220 330578 284226 330580
rect 498193 330578 498259 330581
rect 284220 330576 498259 330578
rect 284220 330520 498198 330576
rect 498254 330520 498259 330576
rect 284220 330518 498259 330520
rect 284220 330516 284226 330518
rect 498193 330515 498259 330518
rect 132493 330442 132559 330445
rect 255814 330442 255820 330444
rect 132493 330440 255820 330442
rect 132493 330384 132498 330440
rect 132554 330384 255820 330440
rect 132493 330382 255820 330384
rect 132493 330379 132559 330382
rect 255814 330380 255820 330382
rect 255884 330380 255890 330444
rect 284702 330380 284708 330444
rect 284772 330442 284778 330444
rect 517513 330442 517579 330445
rect 284772 330440 517579 330442
rect 284772 330384 517518 330440
rect 517574 330384 517579 330440
rect 284772 330382 517579 330384
rect 284772 330380 284778 330382
rect 517513 330379 517579 330382
rect 60825 329218 60891 329221
rect 249517 329218 249583 329221
rect 60825 329216 249583 329218
rect 60825 329160 60830 329216
rect 60886 329160 249522 329216
rect 249578 329160 249583 329216
rect 60825 329158 249583 329160
rect 60825 329155 60891 329158
rect 249517 329155 249583 329158
rect 57973 329082 58039 329085
rect 244733 329082 244799 329085
rect 57973 329080 244799 329082
rect 57973 329024 57978 329080
rect 58034 329024 244738 329080
rect 244794 329024 244799 329080
rect 57973 329022 244799 329024
rect 57973 329019 58039 329022
rect 244733 329019 244799 329022
rect 237373 328266 237439 328269
rect 263910 328266 263916 328268
rect 237373 328264 263916 328266
rect 237373 328208 237378 328264
rect 237434 328208 263916 328264
rect 237373 328206 263916 328208
rect 237373 328203 237439 328206
rect 263910 328204 263916 328206
rect 263980 328204 263986 328268
rect 150433 328130 150499 328133
rect 256918 328130 256924 328132
rect 150433 328128 256924 328130
rect 150433 328072 150438 328128
rect 150494 328072 256924 328128
rect 150433 328070 256924 328072
rect 150433 328067 150499 328070
rect 256918 328068 256924 328070
rect 256988 328068 256994 328132
rect 111793 327994 111859 327997
rect 254894 327994 254900 327996
rect 111793 327992 254900 327994
rect 111793 327936 111798 327992
rect 111854 327936 254900 327992
rect 111793 327934 254900 327936
rect 111793 327931 111859 327934
rect 254894 327932 254900 327934
rect 254964 327932 254970 327996
rect 96613 327858 96679 327861
rect 252870 327858 252876 327860
rect 96613 327856 252876 327858
rect 96613 327800 96618 327856
rect 96674 327800 252876 327856
rect 96613 327798 252876 327800
rect 96613 327795 96679 327798
rect 252870 327796 252876 327798
rect 252940 327796 252946 327860
rect 9673 327722 9739 327725
rect 246246 327722 246252 327724
rect 9673 327720 246252 327722
rect 9673 327664 9678 327720
rect 9734 327664 246252 327720
rect 9673 327662 246252 327664
rect 9673 327659 9739 327662
rect 246246 327660 246252 327662
rect 246316 327660 246322 327724
rect 284886 327660 284892 327724
rect 284956 327722 284962 327724
rect 514753 327722 514819 327725
rect 284956 327720 514819 327722
rect 284956 327664 514758 327720
rect 514814 327664 514819 327720
rect 284956 327662 514819 327664
rect 284956 327660 284962 327662
rect 514753 327659 514819 327662
rect 288709 326770 288775 326773
rect 288709 326768 288818 326770
rect 288709 326712 288714 326768
rect 288770 326712 288818 326768
rect 288709 326707 288818 326712
rect 183553 326634 183619 326637
rect 259862 326634 259868 326636
rect 183553 326632 259868 326634
rect 183553 326576 183558 326632
rect 183614 326576 259868 326632
rect 183553 326574 259868 326576
rect 183553 326571 183619 326574
rect 259862 326572 259868 326574
rect 259932 326572 259938 326636
rect 288758 326501 288818 326707
rect 129733 326498 129799 326501
rect 255630 326498 255636 326500
rect 129733 326496 255636 326498
rect 129733 326440 129738 326496
rect 129794 326440 255636 326496
rect 129733 326438 255636 326440
rect 129733 326435 129799 326438
rect 255630 326436 255636 326438
rect 255700 326436 255706 326500
rect 288709 326496 288818 326501
rect 288709 326440 288714 326496
rect 288770 326440 288818 326496
rect 288709 326438 288818 326440
rect 288709 326435 288775 326438
rect 6913 326362 6979 326365
rect 246062 326362 246068 326364
rect 6913 326360 246068 326362
rect 6913 326304 6918 326360
rect 6974 326304 246068 326360
rect 6913 326302 246068 326304
rect 6913 326299 6979 326302
rect 246062 326300 246068 326302
rect 246132 326300 246138 326364
rect 256049 326362 256115 326365
rect 265566 326362 265572 326364
rect 256049 326360 265572 326362
rect 256049 326304 256054 326360
rect 256110 326304 265572 326360
rect 256049 326302 265572 326304
rect 256049 326299 256115 326302
rect 265566 326300 265572 326302
rect 265636 326300 265642 326364
rect 296621 325820 296687 325821
rect 296621 325818 296668 325820
rect 296576 325816 296668 325818
rect 296732 325818 296738 325820
rect 296576 325760 296626 325816
rect 296576 325758 296668 325760
rect 296621 325756 296668 325758
rect 296732 325758 296814 325818
rect 296732 325756 296738 325758
rect 296621 325755 296687 325756
rect 296621 325682 296687 325685
rect 296576 325680 296730 325682
rect 296576 325624 296626 325680
rect 296682 325624 296730 325680
rect 296576 325622 296730 325624
rect 296621 325619 296730 325622
rect 296670 325548 296730 325619
rect 296662 325484 296668 325548
rect 296732 325484 296738 325548
rect 580257 325274 580323 325277
rect 583520 325274 584960 325364
rect 580257 325272 584960 325274
rect 580257 325216 580262 325272
rect 580318 325216 584960 325272
rect 580257 325214 584960 325216
rect 580257 325211 580323 325214
rect 583520 325124 584960 325214
rect 263501 321604 263567 321605
rect 263501 321602 263548 321604
rect 263456 321600 263548 321602
rect 263456 321544 263506 321600
rect 263456 321542 263548 321544
rect 263501 321540 263548 321542
rect 263612 321540 263618 321604
rect 263501 321539 263567 321540
rect 274030 320724 274036 320788
rect 274100 320786 274106 320788
rect 373993 320786 374059 320789
rect 274100 320784 374059 320786
rect 274100 320728 373998 320784
rect 374054 320728 374059 320784
rect 274100 320726 374059 320728
rect 274100 320724 274106 320726
rect 373993 320723 374059 320726
rect -960 319290 480 319380
rect 3141 319290 3207 319293
rect -960 319288 3207 319290
rect -960 319232 3146 319288
rect 3202 319232 3207 319288
rect -960 319230 3207 319232
rect -960 319140 480 319230
rect 3141 319227 3207 319230
rect 296621 316164 296687 316165
rect 296621 316162 296668 316164
rect 296576 316160 296668 316162
rect 296732 316162 296738 316164
rect 296576 316104 296626 316160
rect 296576 316102 296668 316104
rect 296621 316100 296668 316102
rect 296732 316102 296814 316162
rect 296732 316100 296738 316102
rect 296621 316099 296687 316100
rect 296621 316028 296687 316029
rect 296621 316026 296668 316028
rect 296576 316024 296668 316026
rect 296732 316026 296738 316028
rect 296576 315968 296626 316024
rect 296576 315966 296668 315968
rect 296621 315964 296668 315966
rect 296732 315966 296814 316026
rect 296732 315964 296738 315966
rect 296621 315963 296687 315964
rect 580073 312082 580139 312085
rect 583520 312082 584960 312172
rect 580073 312080 584960 312082
rect 580073 312024 580078 312080
rect 580134 312024 584960 312080
rect 580073 312022 584960 312024
rect 580073 312019 580139 312022
rect 583520 311932 584960 312022
rect 296662 306580 296668 306644
rect 296732 306580 296738 306644
rect 296670 306509 296730 306580
rect 296621 306506 296730 306509
rect 296576 306504 296730 306506
rect 296576 306448 296626 306504
rect 296682 306448 296730 306504
rect 296576 306446 296730 306448
rect 296621 306443 296687 306446
rect 296621 306372 296687 306373
rect 296621 306370 296668 306372
rect 296576 306368 296668 306370
rect 296732 306370 296738 306372
rect -960 306234 480 306324
rect 296576 306312 296626 306368
rect 296576 306310 296668 306312
rect 296621 306308 296668 306310
rect 296732 306310 296814 306370
rect 296732 306308 296738 306310
rect 296621 306307 296687 306308
rect 3325 306234 3391 306237
rect -960 306232 3391 306234
rect -960 306176 3330 306232
rect 3386 306176 3391 306232
rect -960 306174 3391 306176
rect -960 306084 480 306174
rect 3325 306171 3391 306174
rect 580165 298754 580231 298757
rect 583520 298754 584960 298844
rect 580165 298752 584960 298754
rect 580165 298696 580170 298752
rect 580226 298696 584960 298752
rect 580165 298694 584960 298696
rect 580165 298691 580231 298694
rect 583520 298604 584960 298694
rect 296662 296924 296668 296988
rect 296732 296924 296738 296988
rect 296670 296853 296730 296924
rect 296621 296850 296730 296853
rect 296576 296848 296730 296850
rect 296576 296792 296626 296848
rect 296682 296792 296730 296848
rect 296576 296790 296730 296792
rect 296621 296787 296687 296790
rect 296621 296714 296687 296717
rect 296576 296712 296730 296714
rect 296576 296656 296626 296712
rect 296682 296656 296730 296712
rect 296576 296654 296730 296656
rect 296621 296651 296730 296654
rect 296670 296580 296730 296651
rect 296662 296516 296668 296580
rect 296732 296516 296738 296580
rect -960 293178 480 293268
rect 3233 293178 3299 293181
rect -960 293176 3299 293178
rect -960 293120 3238 293176
rect 3294 293120 3299 293176
rect -960 293118 3299 293120
rect -960 293028 480 293118
rect 3233 293115 3299 293118
rect 296621 287196 296687 287197
rect 296621 287194 296668 287196
rect 296576 287192 296668 287194
rect 296732 287194 296738 287196
rect 296576 287136 296626 287192
rect 296576 287134 296668 287136
rect 296621 287132 296668 287134
rect 296732 287134 296814 287194
rect 296732 287132 296738 287134
rect 296621 287131 296687 287132
rect 296621 287058 296687 287061
rect 296576 287056 296730 287058
rect 296576 287000 296626 287056
rect 296682 287000 296730 287056
rect 296576 286998 296730 287000
rect 296621 286995 296730 286998
rect 296670 286924 296730 286995
rect 296662 286860 296668 286924
rect 296732 286860 296738 286924
rect 583520 285276 584960 285516
rect -960 279972 480 280212
rect 296621 277540 296687 277541
rect 296621 277538 296668 277540
rect 296576 277536 296668 277538
rect 296732 277538 296738 277540
rect 296576 277480 296626 277536
rect 296576 277478 296668 277480
rect 296621 277476 296668 277478
rect 296732 277478 296814 277538
rect 296732 277476 296738 277478
rect 296621 277475 296687 277476
rect 296621 277402 296687 277405
rect 296576 277400 296730 277402
rect 296576 277344 296626 277400
rect 296682 277344 296730 277400
rect 296576 277342 296730 277344
rect 296621 277339 296730 277342
rect 296670 277268 296730 277339
rect 296662 277204 296668 277268
rect 296732 277204 296738 277268
rect 580073 272234 580139 272237
rect 583520 272234 584960 272324
rect 580073 272232 584960 272234
rect 580073 272176 580078 272232
rect 580134 272176 584960 272232
rect 580073 272174 584960 272176
rect 580073 272171 580139 272174
rect 583520 272084 584960 272174
rect 296621 267884 296687 267885
rect 296621 267882 296668 267884
rect 296576 267880 296668 267882
rect 296732 267882 296738 267884
rect 296576 267824 296626 267880
rect 296576 267822 296668 267824
rect 296621 267820 296668 267822
rect 296732 267822 296814 267882
rect 296732 267820 296738 267822
rect 296621 267819 296687 267820
rect 296621 267748 296687 267749
rect 296621 267746 296668 267748
rect 296576 267744 296668 267746
rect 296732 267746 296738 267748
rect 296576 267688 296626 267744
rect 296576 267686 296668 267688
rect 296621 267684 296668 267686
rect 296732 267686 296814 267746
rect 296732 267684 296738 267686
rect 296621 267683 296687 267684
rect -960 267202 480 267292
rect 3325 267202 3391 267205
rect -960 267200 3391 267202
rect -960 267144 3330 267200
rect 3386 267144 3391 267200
rect -960 267142 3391 267144
rect -960 267052 480 267142
rect 3325 267139 3391 267142
rect 580073 258906 580139 258909
rect 583520 258906 584960 258996
rect 580073 258904 584960 258906
rect 580073 258848 580078 258904
rect 580134 258848 584960 258904
rect 580073 258846 584960 258848
rect 580073 258843 580139 258846
rect 583520 258756 584960 258846
rect -960 254146 480 254236
rect 3325 254146 3391 254149
rect -960 254144 3391 254146
rect -960 254088 3330 254144
rect 3386 254088 3391 254144
rect -960 254086 3391 254088
rect -960 253996 480 254086
rect 3325 254083 3391 254086
rect 296621 248436 296687 248437
rect 296621 248434 296668 248436
rect 296576 248432 296668 248434
rect 296732 248434 296738 248436
rect 296576 248376 296626 248432
rect 296576 248374 296668 248376
rect 296621 248372 296668 248374
rect 296732 248374 296814 248434
rect 296732 248372 296738 248374
rect 296621 248371 296687 248372
rect 296621 248300 296687 248301
rect 296621 248298 296668 248300
rect 296576 248296 296668 248298
rect 296732 248298 296738 248300
rect 296576 248240 296626 248296
rect 296576 248238 296668 248240
rect 296621 248236 296668 248238
rect 296732 248238 296814 248298
rect 296732 248236 296738 248238
rect 296621 248235 296687 248236
rect 580901 245578 580967 245581
rect 583520 245578 584960 245668
rect 580901 245576 584960 245578
rect 580901 245520 580906 245576
rect 580962 245520 584960 245576
rect 580901 245518 584960 245520
rect 580901 245515 580967 245518
rect 583520 245428 584960 245518
rect -960 241090 480 241180
rect 3325 241090 3391 241093
rect -960 241088 3391 241090
rect -960 241032 3330 241088
rect 3386 241032 3391 241088
rect -960 241030 3391 241032
rect -960 240940 480 241030
rect 3325 241027 3391 241030
rect 296662 238852 296668 238916
rect 296732 238852 296738 238916
rect 296670 238781 296730 238852
rect 296621 238778 296730 238781
rect 296576 238776 296730 238778
rect 296576 238720 296626 238776
rect 296682 238720 296730 238776
rect 296576 238718 296730 238720
rect 296621 238715 296687 238718
rect 296621 238642 296687 238645
rect 296576 238640 296730 238642
rect 296576 238584 296626 238640
rect 296682 238584 296730 238640
rect 296576 238582 296730 238584
rect 296621 238579 296730 238582
rect 296670 238508 296730 238579
rect 296662 238444 296668 238508
rect 296732 238444 296738 238508
rect 580809 232386 580875 232389
rect 583520 232386 584960 232476
rect 580809 232384 584960 232386
rect 580809 232328 580814 232384
rect 580870 232328 584960 232384
rect 580809 232326 584960 232328
rect 580809 232323 580875 232326
rect 583520 232236 584960 232326
rect 296621 229124 296687 229125
rect 296621 229122 296668 229124
rect 296576 229120 296668 229122
rect 296732 229122 296738 229124
rect 296576 229064 296626 229120
rect 296576 229062 296668 229064
rect 296621 229060 296668 229062
rect 296732 229062 296814 229122
rect 296732 229060 296738 229062
rect 296621 229059 296687 229060
rect 296621 228986 296687 228989
rect 296576 228984 296730 228986
rect 296576 228928 296626 228984
rect 296682 228928 296730 228984
rect 296576 228926 296730 228928
rect 296621 228923 296730 228926
rect 296670 228852 296730 228923
rect 296662 228788 296668 228852
rect 296732 228788 296738 228852
rect -960 227884 480 228124
rect 296621 219468 296687 219469
rect 296621 219466 296668 219468
rect 296576 219464 296668 219466
rect 296732 219466 296738 219468
rect 296576 219408 296626 219464
rect 296576 219406 296668 219408
rect 296621 219404 296668 219406
rect 296732 219406 296814 219466
rect 296732 219404 296738 219406
rect 296621 219403 296687 219404
rect 296621 219332 296687 219333
rect 296621 219330 296668 219332
rect 296576 219328 296668 219330
rect 296732 219330 296738 219332
rect 296576 219272 296626 219328
rect 296576 219270 296668 219272
rect 296621 219268 296668 219270
rect 296732 219270 296814 219330
rect 296732 219268 296738 219270
rect 296621 219267 296687 219268
rect 579705 219058 579771 219061
rect 583520 219058 584960 219148
rect 579705 219056 584960 219058
rect 579705 219000 579710 219056
rect 579766 219000 584960 219056
rect 579705 218998 584960 219000
rect 579705 218995 579771 218998
rect 583520 218908 584960 218998
rect -960 214978 480 215068
rect 3325 214978 3391 214981
rect -960 214976 3391 214978
rect -960 214920 3330 214976
rect 3386 214920 3391 214976
rect -960 214918 3391 214920
rect -960 214828 480 214918
rect 3325 214915 3391 214918
rect 237465 214570 237531 214573
rect 238150 214570 238156 214572
rect 237465 214568 238156 214570
rect 237465 214512 237470 214568
rect 237526 214512 238156 214568
rect 237465 214510 238156 214512
rect 237465 214507 237531 214510
rect 238150 214508 238156 214510
rect 238220 214570 238226 214572
rect 335353 214570 335419 214573
rect 238220 214568 335419 214570
rect 238220 214512 335358 214568
rect 335414 214512 335419 214568
rect 238220 214510 335419 214512
rect 238220 214508 238226 214510
rect 335353 214507 335419 214510
rect 296662 209884 296668 209948
rect 296732 209884 296738 209948
rect 296670 209813 296730 209884
rect 296621 209810 296730 209813
rect 296576 209808 296730 209810
rect 296576 209752 296626 209808
rect 296682 209752 296730 209808
rect 296576 209750 296730 209752
rect 296621 209747 296687 209750
rect 296621 209676 296687 209677
rect 296621 209674 296668 209676
rect 296576 209672 296668 209674
rect 296732 209674 296738 209676
rect 296576 209616 296626 209672
rect 296576 209614 296668 209616
rect 296621 209612 296668 209614
rect 296732 209614 296814 209674
rect 296732 209612 296738 209614
rect 296621 209611 296687 209612
rect 580717 205730 580783 205733
rect 583520 205730 584960 205820
rect 580717 205728 584960 205730
rect 580717 205672 580722 205728
rect 580778 205672 584960 205728
rect 580717 205670 584960 205672
rect 580717 205667 580783 205670
rect 583520 205580 584960 205670
rect -960 201922 480 202012
rect 3693 201922 3759 201925
rect -960 201920 3759 201922
rect -960 201864 3698 201920
rect 3754 201864 3759 201920
rect -960 201862 3759 201864
rect -960 201772 480 201862
rect 3693 201859 3759 201862
rect 296662 200228 296668 200292
rect 296732 200228 296738 200292
rect 296670 200157 296730 200228
rect 296621 200154 296730 200157
rect 296576 200152 296730 200154
rect 296576 200096 296626 200152
rect 296682 200096 296730 200152
rect 296576 200094 296730 200096
rect 296621 200091 296687 200094
rect 296621 200020 296687 200021
rect 296621 200018 296668 200020
rect 296576 200016 296668 200018
rect 296732 200018 296738 200020
rect 296576 199960 296626 200016
rect 296576 199958 296668 199960
rect 296621 199956 296668 199958
rect 296732 199958 296814 200018
rect 296732 199956 296738 199958
rect 296621 199955 296687 199956
rect 287697 194578 287763 194581
rect 293902 194578 293908 194580
rect 287697 194576 293908 194578
rect 287697 194520 287702 194576
rect 287758 194520 293908 194576
rect 287697 194518 293908 194520
rect 287697 194515 287763 194518
rect 293902 194516 293908 194518
rect 293972 194516 293978 194580
rect 580533 192538 580599 192541
rect 583520 192538 584960 192628
rect 580533 192536 584960 192538
rect 580533 192480 580538 192536
rect 580594 192480 584960 192536
rect 580533 192478 584960 192480
rect 580533 192475 580599 192478
rect 583520 192388 584960 192478
rect 296662 190572 296668 190636
rect 296732 190572 296738 190636
rect 296670 190501 296730 190572
rect 296621 190498 296730 190501
rect 296576 190496 296730 190498
rect 296576 190440 296626 190496
rect 296682 190440 296730 190496
rect 296576 190438 296730 190440
rect 296621 190435 296687 190438
rect 296621 190362 296687 190365
rect 296576 190360 296730 190362
rect 296576 190304 296626 190360
rect 296682 190304 296730 190360
rect 296576 190302 296730 190304
rect 296621 190299 296730 190302
rect 296670 190228 296730 190299
rect 296662 190164 296668 190228
rect 296732 190164 296738 190228
rect -960 188866 480 188956
rect 3601 188866 3667 188869
rect -960 188864 3667 188866
rect -960 188808 3606 188864
rect 3662 188808 3667 188864
rect -960 188806 3667 188808
rect -960 188716 480 188806
rect 3601 188803 3667 188806
rect 279734 186900 279740 186964
rect 279804 186962 279810 186964
rect 444373 186962 444439 186965
rect 279804 186960 444439 186962
rect 279804 186904 444378 186960
rect 444434 186904 444439 186960
rect 279804 186902 444439 186904
rect 279804 186900 279810 186902
rect 444373 186899 444439 186902
rect 296621 180844 296687 180845
rect 296621 180842 296668 180844
rect 296576 180840 296668 180842
rect 296732 180842 296738 180844
rect 296576 180784 296626 180840
rect 296576 180782 296668 180784
rect 296621 180780 296668 180782
rect 296732 180782 296814 180842
rect 296732 180780 296738 180782
rect 296621 180779 296687 180780
rect 296621 180706 296687 180709
rect 296576 180704 296730 180706
rect 296576 180648 296626 180704
rect 296682 180648 296730 180704
rect 296576 180646 296730 180648
rect 296621 180643 296730 180646
rect 296670 180572 296730 180643
rect 296662 180508 296668 180572
rect 296732 180508 296738 180572
rect 293350 179964 293356 180028
rect 293420 180026 293426 180028
rect 345381 180026 345447 180029
rect 293420 180024 345447 180026
rect 293420 179968 345386 180024
rect 345442 179968 345447 180024
rect 293420 179966 345447 179968
rect 293420 179964 293426 179966
rect 345381 179963 345447 179966
rect 579705 179210 579771 179213
rect 583520 179210 584960 179300
rect 579705 179208 584960 179210
rect 579705 179152 579710 179208
rect 579766 179152 584960 179208
rect 579705 179150 584960 179152
rect 579705 179147 579771 179150
rect 583520 179060 584960 179150
rect 62113 177306 62179 177309
rect 250294 177306 250300 177308
rect 62113 177304 250300 177306
rect 62113 177248 62118 177304
rect 62174 177248 250300 177304
rect 62113 177246 250300 177248
rect 62113 177243 62179 177246
rect 250294 177244 250300 177246
rect 250364 177244 250370 177308
rect 288014 177244 288020 177308
rect 288084 177306 288090 177308
rect 553393 177306 553459 177309
rect 288084 177304 553459 177306
rect 288084 177248 553398 177304
rect 553454 177248 553459 177304
rect 288084 177246 553459 177248
rect 288084 177244 288090 177246
rect 553393 177243 553459 177246
rect -960 175796 480 176036
rect 276054 175884 276060 175948
rect 276124 175946 276130 175948
rect 407205 175946 407271 175949
rect 276124 175944 407271 175946
rect 276124 175888 407210 175944
rect 407266 175888 407271 175944
rect 276124 175886 407271 175888
rect 276124 175884 276130 175886
rect 407205 175883 407271 175886
rect 274214 174660 274220 174724
rect 274284 174722 274290 174724
rect 374085 174722 374151 174725
rect 274284 174720 374151 174722
rect 274284 174664 374090 174720
rect 374146 174664 374151 174720
rect 274284 174662 374151 174664
rect 274284 174660 274290 174662
rect 374085 174659 374151 174662
rect 283782 174524 283788 174588
rect 283852 174586 283858 174588
rect 499573 174586 499639 174589
rect 283852 174584 499639 174586
rect 283852 174528 499578 174584
rect 499634 174528 499639 174584
rect 283852 174526 499639 174528
rect 283852 174524 283858 174526
rect 499573 174523 499639 174526
rect 283966 173436 283972 173500
rect 284036 173498 284042 173500
rect 496813 173498 496879 173501
rect 284036 173496 496879 173498
rect 284036 173440 496818 173496
rect 496874 173440 496879 173496
rect 284036 173438 496879 173440
rect 284036 173436 284042 173438
rect 496813 173435 496879 173438
rect 286174 173300 286180 173364
rect 286244 173362 286250 173364
rect 534073 173362 534139 173365
rect 286244 173360 534139 173362
rect 286244 173304 534078 173360
rect 534134 173304 534139 173360
rect 286244 173302 534139 173304
rect 286244 173300 286250 173302
rect 534073 173299 534139 173302
rect 289302 173164 289308 173228
rect 289372 173226 289378 173228
rect 569953 173226 570019 173229
rect 289372 173224 570019 173226
rect 289372 173168 569958 173224
rect 570014 173168 570019 173224
rect 289372 173166 570019 173168
rect 289372 173164 289378 173166
rect 569953 173163 570019 173166
rect 296621 171188 296687 171189
rect 296621 171186 296668 171188
rect 296576 171184 296668 171186
rect 296732 171186 296738 171188
rect 296576 171128 296626 171184
rect 296576 171126 296668 171128
rect 296621 171124 296668 171126
rect 296732 171126 296814 171186
rect 296732 171124 296738 171126
rect 296621 171123 296687 171124
rect 296621 171052 296687 171053
rect 296621 171050 296668 171052
rect 296576 171048 296668 171050
rect 296732 171050 296738 171052
rect 296576 170992 296626 171048
rect 296576 170990 296668 170992
rect 296621 170988 296668 170990
rect 296732 170990 296814 171050
rect 296732 170988 296738 170990
rect 296621 170987 296687 170988
rect 295006 170444 295012 170508
rect 295076 170506 295082 170508
rect 345473 170506 345539 170509
rect 295076 170504 345539 170506
rect 295076 170448 345478 170504
rect 345534 170448 345539 170504
rect 295076 170446 345539 170448
rect 295076 170444 295082 170446
rect 345473 170443 345539 170446
rect 282494 170308 282500 170372
rect 282564 170370 282570 170372
rect 481633 170370 481699 170373
rect 282564 170368 481699 170370
rect 282564 170312 481638 170368
rect 481694 170312 481699 170368
rect 282564 170310 481699 170312
rect 282564 170308 282570 170310
rect 481633 170307 481699 170310
rect 278446 166500 278452 166564
rect 278516 166562 278522 166564
rect 425053 166562 425119 166565
rect 278516 166560 425119 166562
rect 278516 166504 425058 166560
rect 425114 166504 425119 166560
rect 278516 166502 425119 166504
rect 278516 166500 278522 166502
rect 425053 166499 425119 166502
rect 278630 166364 278636 166428
rect 278700 166426 278706 166428
rect 426433 166426 426499 166429
rect 278700 166424 426499 166426
rect 278700 166368 426438 166424
rect 426494 166368 426499 166424
rect 278700 166366 426499 166368
rect 278700 166364 278706 166366
rect 426433 166363 426499 166366
rect 279550 166228 279556 166292
rect 279620 166290 279626 166292
rect 447133 166290 447199 166293
rect 279620 166288 447199 166290
rect 279620 166232 447138 166288
rect 447194 166232 447199 166288
rect 279620 166230 447199 166232
rect 279620 166228 279626 166230
rect 447133 166227 447199 166230
rect 580165 165882 580231 165885
rect 583520 165882 584960 165972
rect 580165 165880 584960 165882
rect 580165 165824 580170 165880
rect 580226 165824 584960 165880
rect 580165 165822 584960 165824
rect 580165 165819 580231 165822
rect 583520 165732 584960 165822
rect 274398 165004 274404 165068
rect 274468 165066 274474 165068
rect 375373 165066 375439 165069
rect 274468 165064 375439 165066
rect 274468 165008 375378 165064
rect 375434 165008 375439 165064
rect 274468 165006 375439 165008
rect 274468 165004 274474 165006
rect 375373 165003 375439 165006
rect 275870 164868 275876 164932
rect 275940 164930 275946 164932
rect 390553 164930 390619 164933
rect 275940 164928 390619 164930
rect 275940 164872 390558 164928
rect 390614 164872 390619 164928
rect 275940 164870 390619 164872
rect 275940 164868 275946 164870
rect 390553 164867 390619 164870
rect 257337 163434 257403 163437
rect 296846 163434 296852 163436
rect 257337 163432 296852 163434
rect 257337 163376 257342 163432
rect 257398 163376 296852 163432
rect 257337 163374 296852 163376
rect 257337 163371 257403 163374
rect 296846 163372 296852 163374
rect 296916 163372 296922 163436
rect -960 162890 480 162980
rect 3325 162890 3391 162893
rect -960 162888 3391 162890
rect -960 162832 3330 162888
rect 3386 162832 3391 162888
rect -960 162830 3391 162832
rect -960 162740 480 162830
rect 3325 162827 3391 162830
rect 285070 162284 285076 162348
rect 285140 162346 285146 162348
rect 514845 162346 514911 162349
rect 285140 162344 514911 162346
rect 285140 162288 514850 162344
rect 514906 162288 514911 162344
rect 285140 162286 514911 162288
rect 285140 162284 285146 162286
rect 514845 162283 514911 162286
rect 286726 162148 286732 162212
rect 286796 162210 286802 162212
rect 531405 162210 531471 162213
rect 286796 162208 531471 162210
rect 286796 162152 531410 162208
rect 531466 162152 531471 162208
rect 286796 162150 531471 162152
rect 286796 162148 286802 162150
rect 531405 162147 531471 162150
rect 289486 162012 289492 162076
rect 289556 162074 289562 162076
rect 568573 162074 568639 162077
rect 289556 162072 568639 162074
rect 289556 162016 568578 162072
rect 568634 162016 568639 162072
rect 289556 162014 568639 162016
rect 289556 162012 289562 162014
rect 568573 162011 568639 162014
rect 296621 161530 296687 161533
rect 296846 161530 296852 161532
rect 296576 161528 296852 161530
rect 296576 161472 296626 161528
rect 296682 161472 296852 161528
rect 296576 161470 296852 161472
rect 296621 161467 296687 161470
rect 296846 161468 296852 161470
rect 296916 161468 296922 161532
rect 241145 161394 241211 161397
rect 269573 161394 269639 161397
rect 241145 161392 269639 161394
rect 241145 161336 241150 161392
rect 241206 161336 269578 161392
rect 269634 161336 269639 161392
rect 241145 161334 269639 161336
rect 241145 161331 241211 161334
rect 269573 161331 269639 161334
rect 296110 161332 296116 161396
rect 296180 161394 296186 161396
rect 296478 161394 296484 161396
rect 296180 161334 296484 161394
rect 296180 161332 296186 161334
rect 296478 161332 296484 161334
rect 296548 161332 296554 161396
rect 301773 161394 301839 161397
rect 345422 161394 345428 161396
rect 301773 161392 345428 161394
rect 301773 161336 301778 161392
rect 301834 161336 345428 161392
rect 301773 161334 345428 161336
rect 301773 161331 301839 161334
rect 345422 161332 345428 161334
rect 345492 161332 345498 161396
rect 241237 161258 241303 161261
rect 269849 161258 269915 161261
rect 241237 161256 269915 161258
rect 241237 161200 241242 161256
rect 241298 161200 269854 161256
rect 269910 161200 269915 161256
rect 241237 161198 269915 161200
rect 241237 161195 241303 161198
rect 269849 161195 269915 161198
rect 290958 161196 290964 161260
rect 291028 161258 291034 161260
rect 348325 161258 348391 161261
rect 291028 161256 348391 161258
rect 291028 161200 348330 161256
rect 348386 161200 348391 161256
rect 291028 161198 348391 161200
rect 291028 161196 291034 161198
rect 348325 161195 348391 161198
rect 239581 161122 239647 161125
rect 268510 161122 268516 161124
rect 239581 161120 268516 161122
rect 239581 161064 239586 161120
rect 239642 161064 268516 161120
rect 239581 161062 268516 161064
rect 239581 161059 239647 161062
rect 268510 161060 268516 161062
rect 268580 161060 268586 161124
rect 272333 161122 272399 161125
rect 343582 161122 343588 161124
rect 272333 161120 343588 161122
rect 272333 161064 272338 161120
rect 272394 161064 343588 161120
rect 272333 161062 343588 161064
rect 272333 161059 272399 161062
rect 343582 161060 343588 161062
rect 343652 161060 343658 161124
rect 262622 160924 262628 160988
rect 262692 160986 262698 160988
rect 349429 160986 349495 160989
rect 262692 160984 349495 160986
rect 262692 160928 349434 160984
rect 349490 160928 349495 160984
rect 262692 160926 349495 160928
rect 262692 160924 262698 160926
rect 349429 160923 349495 160926
rect 239857 160850 239923 160853
rect 269665 160850 269731 160853
rect 239857 160848 269731 160850
rect 239857 160792 239862 160848
rect 239918 160792 269670 160848
rect 269726 160792 269731 160848
rect 239857 160790 269731 160792
rect 239857 160787 239923 160790
rect 269665 160787 269731 160790
rect 282678 160788 282684 160852
rect 282748 160850 282754 160852
rect 481725 160850 481791 160853
rect 282748 160848 481791 160850
rect 282748 160792 481730 160848
rect 481786 160792 481791 160848
rect 282748 160790 481791 160792
rect 282748 160788 282754 160790
rect 481725 160787 481791 160790
rect 215293 160714 215359 160717
rect 261385 160714 261451 160717
rect 215293 160712 261451 160714
rect 215293 160656 215298 160712
rect 215354 160656 261390 160712
rect 261446 160656 261451 160712
rect 215293 160654 261451 160656
rect 215293 160651 215359 160654
rect 261385 160651 261451 160654
rect 287830 160652 287836 160716
rect 287900 160714 287906 160716
rect 550633 160714 550699 160717
rect 287900 160712 550699 160714
rect 287900 160656 550638 160712
rect 550694 160656 550699 160712
rect 287900 160654 550699 160656
rect 287900 160652 287906 160654
rect 550633 160651 550699 160654
rect 245561 160578 245627 160581
rect 269757 160578 269823 160581
rect 245561 160576 269823 160578
rect 245561 160520 245566 160576
rect 245622 160520 269762 160576
rect 269818 160520 269823 160576
rect 245561 160518 269823 160520
rect 245561 160515 245627 160518
rect 269757 160515 269823 160518
rect 277158 159564 277164 159628
rect 277228 159626 277234 159628
rect 409873 159626 409939 159629
rect 277228 159624 409939 159626
rect 277228 159568 409878 159624
rect 409934 159568 409939 159624
rect 277228 159566 409939 159568
rect 277228 159564 277234 159566
rect 409873 159563 409939 159566
rect 255681 159490 255747 159493
rect 265198 159490 265204 159492
rect 255681 159488 265204 159490
rect 255681 159432 255686 159488
rect 255742 159432 265204 159488
rect 255681 159430 265204 159432
rect 255681 159427 255747 159430
rect 265198 159428 265204 159430
rect 265268 159428 265274 159492
rect 286910 159428 286916 159492
rect 286980 159490 286986 159492
rect 532693 159490 532759 159493
rect 286980 159488 532759 159490
rect 286980 159432 532698 159488
rect 532754 159432 532759 159488
rect 286980 159430 532759 159432
rect 286980 159428 286986 159430
rect 532693 159427 532759 159430
rect 235993 159354 236059 159357
rect 263726 159354 263732 159356
rect 235993 159352 263732 159354
rect 235993 159296 235998 159352
rect 236054 159296 263732 159352
rect 235993 159294 263732 159296
rect 235993 159291 236059 159294
rect 263726 159292 263732 159294
rect 263796 159292 263802 159356
rect 296294 159292 296300 159356
rect 296364 159354 296370 159356
rect 580533 159354 580599 159357
rect 296364 159352 580599 159354
rect 296364 159296 580538 159352
rect 580594 159296 580599 159352
rect 296364 159294 580599 159296
rect 296364 159292 296370 159294
rect 580533 159291 580599 159294
rect 258441 158810 258507 158813
rect 265382 158810 265388 158812
rect 258441 158808 265388 158810
rect 258441 158752 258446 158808
rect 258502 158752 265388 158808
rect 258441 158750 265388 158752
rect 258441 158747 258507 158750
rect 265382 158748 265388 158750
rect 265452 158748 265458 158812
rect 253105 158674 253171 158677
rect 265014 158674 265020 158676
rect 253105 158672 265020 158674
rect 253105 158616 253110 158672
rect 253166 158616 265020 158672
rect 253105 158614 265020 158616
rect 253105 158611 253171 158614
rect 265014 158612 265020 158614
rect 265084 158612 265090 158676
rect 269021 158674 269087 158677
rect 295742 158674 295748 158676
rect 269021 158672 295748 158674
rect 269021 158616 269026 158672
rect 269082 158616 295748 158672
rect 269021 158614 295748 158616
rect 269021 158611 269087 158614
rect 295742 158612 295748 158614
rect 295812 158612 295818 158676
rect 296662 158612 296668 158676
rect 296732 158674 296738 158676
rect 298001 158674 298067 158677
rect 296732 158672 298067 158674
rect 296732 158616 298006 158672
rect 298062 158616 298067 158672
rect 296732 158614 298067 158616
rect 296732 158612 296738 158614
rect 298001 158611 298067 158614
rect 258993 158538 259059 158541
rect 291142 158538 291148 158540
rect 258993 158536 291148 158538
rect 258993 158480 258998 158536
rect 259054 158480 291148 158536
rect 258993 158478 291148 158480
rect 258993 158475 259059 158478
rect 291142 158476 291148 158478
rect 291212 158476 291218 158540
rect 293166 158476 293172 158540
rect 293236 158538 293242 158540
rect 310881 158538 310947 158541
rect 293236 158536 310947 158538
rect 293236 158480 310886 158536
rect 310942 158480 310947 158536
rect 293236 158478 310947 158480
rect 293236 158476 293242 158478
rect 310881 158475 310947 158478
rect 234061 158402 234127 158405
rect 277393 158402 277459 158405
rect 234061 158400 277459 158402
rect 234061 158344 234066 158400
rect 234122 158344 277398 158400
rect 277454 158344 277459 158400
rect 234061 158342 277459 158344
rect 234061 158339 234127 158342
rect 277393 158339 277459 158342
rect 288750 158340 288756 158404
rect 288820 158402 288826 158404
rect 289629 158402 289695 158405
rect 288820 158400 289695 158402
rect 288820 158344 289634 158400
rect 289690 158344 289695 158400
rect 288820 158342 289695 158344
rect 288820 158340 288826 158342
rect 289629 158339 289695 158342
rect 290590 158340 290596 158404
rect 290660 158402 290666 158404
rect 343633 158402 343699 158405
rect 290660 158400 343699 158402
rect 290660 158344 343638 158400
rect 343694 158344 343699 158400
rect 290660 158342 343699 158344
rect 290660 158340 290666 158342
rect 343633 158339 343699 158342
rect 248321 158266 248387 158269
rect 266486 158266 266492 158268
rect 248321 158264 266492 158266
rect 248321 158208 248326 158264
rect 248382 158208 266492 158264
rect 248321 158206 266492 158208
rect 248321 158203 248387 158206
rect 266486 158204 266492 158206
rect 266556 158204 266562 158268
rect 271638 158204 271644 158268
rect 271708 158266 271714 158268
rect 345289 158266 345355 158269
rect 271708 158264 345355 158266
rect 271708 158208 345294 158264
rect 345350 158208 345355 158264
rect 271708 158206 345355 158208
rect 271708 158204 271714 158206
rect 345289 158203 345355 158206
rect 238753 158130 238819 158133
rect 263542 158130 263548 158132
rect 238753 158128 263548 158130
rect 238753 158072 238758 158128
rect 238814 158072 263548 158128
rect 238753 158070 263548 158072
rect 238753 158067 238819 158070
rect 263542 158068 263548 158070
rect 263612 158068 263618 158132
rect 270166 158068 270172 158132
rect 270236 158130 270242 158132
rect 348141 158130 348207 158133
rect 270236 158128 348207 158130
rect 270236 158072 348146 158128
rect 348202 158072 348207 158128
rect 270236 158070 348207 158072
rect 270236 158068 270242 158070
rect 348141 158067 348207 158070
rect 218145 157994 218211 157997
rect 262254 157994 262260 157996
rect 218145 157992 262260 157994
rect 218145 157936 218150 157992
rect 218206 157936 262260 157992
rect 218145 157934 262260 157936
rect 218145 157931 218211 157934
rect 262254 157932 262260 157934
rect 262324 157932 262330 157996
rect 284385 157994 284451 157997
rect 507853 157994 507919 157997
rect 284385 157992 507919 157994
rect 284385 157936 284390 157992
rect 284446 157936 507858 157992
rect 507914 157936 507919 157992
rect 284385 157934 507919 157936
rect 284385 157931 284451 157934
rect 507853 157931 507919 157934
rect 291694 157796 291700 157860
rect 291764 157858 291770 157860
rect 302509 157858 302575 157861
rect 291764 157856 302575 157858
rect 291764 157800 302514 157856
rect 302570 157800 302575 157856
rect 291764 157798 302575 157800
rect 291764 157796 291770 157798
rect 302509 157795 302575 157798
rect 343725 157450 343791 157453
rect 344686 157450 344692 157452
rect 343725 157448 344692 157450
rect 343725 157392 343730 157448
rect 343786 157392 344692 157448
rect 343725 157390 344692 157392
rect 343725 157387 343791 157390
rect 344686 157388 344692 157390
rect 344756 157388 344762 157452
rect 201493 156634 201559 156637
rect 260966 156634 260972 156636
rect 201493 156632 260972 156634
rect 201493 156576 201498 156632
rect 201554 156576 260972 156632
rect 201493 156574 260972 156576
rect 201493 156571 201559 156574
rect 260966 156572 260972 156574
rect 261036 156572 261042 156636
rect 283598 156572 283604 156636
rect 283668 156634 283674 156636
rect 498285 156634 498351 156637
rect 283668 156632 498351 156634
rect 283668 156576 498290 156632
rect 498346 156576 498351 156632
rect 283668 156574 498351 156576
rect 283668 156572 283674 156574
rect 498285 156571 498351 156574
rect 257429 155954 257495 155957
rect 268326 155954 268332 155956
rect 257429 155952 268332 155954
rect 257429 155896 257434 155952
rect 257490 155896 268332 155952
rect 257429 155894 268332 155896
rect 257429 155891 257495 155894
rect 268326 155892 268332 155894
rect 268396 155892 268402 155956
rect 257838 155756 257844 155820
rect 257908 155818 257914 155820
rect 269297 155818 269363 155821
rect 257908 155816 269363 155818
rect 257908 155760 269302 155816
rect 269358 155760 269363 155816
rect 257908 155758 269363 155760
rect 257908 155756 257914 155758
rect 269297 155755 269363 155758
rect 209865 155682 209931 155685
rect 260281 155682 260347 155685
rect 209865 155680 260347 155682
rect 209865 155624 209870 155680
rect 209926 155624 260286 155680
rect 260342 155624 260347 155680
rect 209865 155622 260347 155624
rect 209865 155619 209931 155622
rect 260281 155619 260347 155622
rect 260414 155620 260420 155684
rect 260484 155682 260490 155684
rect 266445 155682 266511 155685
rect 260484 155680 266511 155682
rect 260484 155624 266450 155680
rect 266506 155624 266511 155680
rect 260484 155622 266511 155624
rect 260484 155620 260490 155622
rect 266445 155619 266511 155622
rect 284017 155682 284083 155685
rect 284150 155682 284156 155684
rect 284017 155680 284156 155682
rect 284017 155624 284022 155680
rect 284078 155624 284156 155680
rect 284017 155622 284156 155624
rect 284017 155619 284083 155622
rect 284150 155620 284156 155622
rect 284220 155620 284226 155684
rect 296110 155620 296116 155684
rect 296180 155682 296186 155684
rect 349889 155682 349955 155685
rect 296180 155680 349955 155682
rect 296180 155624 349894 155680
rect 349950 155624 349955 155680
rect 296180 155622 349955 155624
rect 296180 155620 296186 155622
rect 349889 155619 349955 155622
rect 201585 155546 201651 155549
rect 261150 155546 261156 155548
rect 201585 155544 261156 155546
rect 201585 155488 201590 155544
rect 201646 155488 261156 155544
rect 201585 155486 261156 155488
rect 201585 155483 201651 155486
rect 261150 155484 261156 155486
rect 261220 155484 261226 155548
rect 270350 155484 270356 155548
rect 270420 155546 270426 155548
rect 345841 155546 345907 155549
rect 270420 155544 345907 155546
rect 270420 155488 345846 155544
rect 345902 155488 345907 155544
rect 270420 155486 345907 155488
rect 270420 155484 270426 155486
rect 345841 155483 345907 155486
rect 186313 155410 186379 155413
rect 259678 155410 259684 155412
rect 186313 155408 259684 155410
rect 186313 155352 186318 155408
rect 186374 155352 259684 155408
rect 186313 155350 259684 155352
rect 186313 155347 186379 155350
rect 259678 155348 259684 155350
rect 259748 155348 259754 155412
rect 260598 155348 260604 155412
rect 260668 155410 260674 155412
rect 269389 155410 269455 155413
rect 260668 155408 269455 155410
rect 260668 155352 269394 155408
rect 269450 155352 269455 155408
rect 260668 155350 269455 155352
rect 260668 155348 260674 155350
rect 269389 155347 269455 155350
rect 273161 155410 273227 155413
rect 356053 155410 356119 155413
rect 273161 155408 356119 155410
rect 273161 155352 273166 155408
rect 273222 155352 356058 155408
rect 356114 155352 356119 155408
rect 273161 155350 356119 155352
rect 273161 155347 273227 155350
rect 356053 155347 356119 155350
rect 185025 155274 185091 155277
rect 259494 155274 259500 155276
rect 185025 155272 259500 155274
rect 185025 155216 185030 155272
rect 185086 155216 259500 155272
rect 185025 155214 259500 155216
rect 185025 155211 185091 155214
rect 259494 155212 259500 155214
rect 259564 155212 259570 155276
rect 284150 155212 284156 155276
rect 284220 155274 284226 155276
rect 494053 155274 494119 155277
rect 284220 155272 494119 155274
rect 284220 155216 494058 155272
rect 494114 155216 494119 155272
rect 284220 155214 494119 155216
rect 284220 155212 284226 155214
rect 494053 155211 494119 155214
rect 257613 155138 257679 155141
rect 266302 155138 266308 155140
rect 257613 155136 266308 155138
rect 257613 155080 257618 155136
rect 257674 155080 266308 155136
rect 257613 155078 266308 155080
rect 257613 155075 257679 155078
rect 266302 155076 266308 155078
rect 266372 155076 266378 155140
rect 257654 153852 257660 153916
rect 257724 153914 257730 153916
rect 269062 153914 269068 153916
rect 257724 153854 269068 153914
rect 257724 153852 257730 153854
rect 269062 153852 269068 153854
rect 269132 153852 269138 153916
rect 248229 153778 248295 153781
rect 268142 153778 268148 153780
rect 248229 153776 268148 153778
rect 248229 153720 248234 153776
rect 248290 153720 268148 153776
rect 248229 153718 268148 153720
rect 248229 153715 248295 153718
rect 268142 153716 268148 153718
rect 268212 153716 268218 153780
rect 580625 152690 580691 152693
rect 583520 152690 584960 152780
rect 580625 152688 584960 152690
rect 580625 152632 580630 152688
rect 580686 152632 584960 152688
rect 580625 152630 584960 152632
rect 580625 152627 580691 152630
rect 583520 152540 584960 152630
rect 256693 152418 256759 152421
rect 256693 152416 260084 152418
rect 256693 152360 256698 152416
rect 256754 152360 260084 152416
rect 256693 152358 260084 152360
rect 256693 152355 256759 152358
rect 257470 151812 257476 151876
rect 257540 151874 257546 151876
rect 258022 151874 258028 151876
rect 257540 151814 258028 151874
rect 257540 151812 257546 151814
rect 258022 151812 258028 151814
rect 258092 151812 258098 151876
rect 257470 151676 257476 151740
rect 257540 151738 257546 151740
rect 258022 151738 258028 151740
rect 257540 151678 258028 151738
rect 257540 151676 257546 151678
rect 258022 151676 258028 151678
rect 258092 151676 258098 151740
rect 344645 151738 344711 151741
rect 343804 151736 344711 151738
rect 343804 151680 344650 151736
rect 344706 151680 344711 151736
rect 343804 151678 344711 151680
rect 344645 151675 344711 151678
rect -960 149834 480 149924
rect 3325 149834 3391 149837
rect -960 149832 3391 149834
rect -960 149776 3330 149832
rect 3386 149776 3391 149832
rect -960 149774 3391 149776
rect -960 149684 480 149774
rect 3325 149771 3391 149774
rect 257245 148338 257311 148341
rect 257245 148336 260084 148338
rect 257245 148280 257250 148336
rect 257306 148280 260084 148336
rect 257245 148278 260084 148280
rect 257245 148275 257311 148278
rect 343398 148276 343404 148340
rect 343468 148338 343474 148340
rect 344645 148338 344711 148341
rect 343468 148336 344711 148338
rect 343468 148280 344650 148336
rect 344706 148280 344711 148336
rect 343468 148278 344711 148280
rect 343468 148276 343474 148278
rect 344645 148275 344711 148278
rect 345105 147658 345171 147661
rect 343804 147656 345171 147658
rect 343804 147600 345110 147656
rect 345166 147600 345171 147656
rect 343804 147598 345171 147600
rect 345105 147595 345171 147598
rect 256693 143578 256759 143581
rect 256693 143576 260084 143578
rect 256693 143520 256698 143576
rect 256754 143520 260084 143576
rect 256693 143518 260084 143520
rect 256693 143515 256759 143518
rect 345238 142898 345244 142900
rect 343804 142838 345244 142898
rect 345238 142836 345244 142838
rect 345308 142836 345314 142900
rect 257470 142156 257476 142220
rect 257540 142218 257546 142220
rect 258022 142218 258028 142220
rect 257540 142158 258028 142218
rect 257540 142156 257546 142158
rect 258022 142156 258028 142158
rect 258092 142156 258098 142220
rect 257797 141946 257863 141949
rect 258022 141946 258028 141948
rect 257797 141944 258028 141946
rect 257797 141888 257802 141944
rect 257858 141888 258028 141944
rect 257797 141886 258028 141888
rect 257797 141883 257863 141886
rect 258022 141884 258028 141886
rect 258092 141884 258098 141948
rect 257245 139498 257311 139501
rect 257245 139496 260084 139498
rect 257245 139440 257250 139496
rect 257306 139440 260084 139496
rect 257245 139438 260084 139440
rect 257245 139435 257311 139438
rect 579613 139362 579679 139365
rect 583520 139362 584960 139452
rect 579613 139360 584960 139362
rect 579613 139304 579618 139360
rect 579674 139304 584960 139360
rect 579613 139302 584960 139304
rect 579613 139299 579679 139302
rect 583520 139212 584960 139302
rect 345749 138818 345815 138821
rect 343804 138816 345815 138818
rect 343804 138760 345754 138816
rect 345810 138760 345815 138816
rect 343804 138758 345815 138760
rect 345749 138755 345815 138758
rect -960 136778 480 136868
rect 3049 136778 3115 136781
rect -960 136776 3115 136778
rect -960 136720 3054 136776
rect 3110 136720 3115 136776
rect -960 136718 3115 136720
rect -960 136628 480 136718
rect 3049 136715 3115 136718
rect 256785 134738 256851 134741
rect 256785 134736 260084 134738
rect 256785 134680 256790 134736
rect 256846 134680 260084 134736
rect 256785 134678 260084 134680
rect 256785 134675 256851 134678
rect 345013 134058 345079 134061
rect 343804 134056 345079 134058
rect 343804 134000 345018 134056
rect 345074 134000 345079 134056
rect 343804 133998 345079 134000
rect 345013 133995 345079 133998
rect 257797 132562 257863 132565
rect 258022 132562 258028 132564
rect 257797 132560 258028 132562
rect 257797 132504 257802 132560
rect 257858 132504 258028 132560
rect 257797 132502 258028 132504
rect 257797 132499 257863 132502
rect 258022 132500 258028 132502
rect 258092 132500 258098 132564
rect 257797 132426 257863 132429
rect 258022 132426 258028 132428
rect 257797 132424 258028 132426
rect 257797 132368 257802 132424
rect 257858 132368 258028 132424
rect 257797 132366 258028 132368
rect 257797 132363 257863 132366
rect 258022 132364 258028 132366
rect 258092 132364 258098 132428
rect 256785 130658 256851 130661
rect 256785 130656 260084 130658
rect 256785 130600 256790 130656
rect 256846 130600 260084 130656
rect 256785 130598 260084 130600
rect 256785 130595 256851 130598
rect 345565 129978 345631 129981
rect 343804 129976 345631 129978
rect 343804 129920 345570 129976
rect 345626 129920 345631 129976
rect 343804 129918 345631 129920
rect 345565 129915 345631 129918
rect 344686 129780 344692 129844
rect 344756 129842 344762 129844
rect 344921 129842 344987 129845
rect 344756 129840 344987 129842
rect 344756 129784 344926 129840
rect 344982 129784 344987 129840
rect 344756 129782 344987 129784
rect 344756 129780 344762 129782
rect 344921 129779 344987 129782
rect 579705 126034 579771 126037
rect 583520 126034 584960 126124
rect 579705 126032 584960 126034
rect 579705 125976 579710 126032
rect 579766 125976 584960 126032
rect 579705 125974 584960 125976
rect 579705 125971 579771 125974
rect 256785 125898 256851 125901
rect 256785 125896 260084 125898
rect 256785 125840 256790 125896
rect 256846 125840 260084 125896
rect 583520 125884 584960 125974
rect 256785 125838 260084 125840
rect 256785 125835 256851 125838
rect 345473 125218 345539 125221
rect 343804 125216 345539 125218
rect 343804 125160 345478 125216
rect 345534 125160 345539 125216
rect 343804 125158 345539 125160
rect 345473 125155 345539 125158
rect -960 123572 480 123812
rect 257797 122906 257863 122909
rect 258022 122906 258028 122908
rect 257797 122904 258028 122906
rect 257797 122848 257802 122904
rect 257858 122848 258028 122904
rect 257797 122846 258028 122848
rect 257797 122843 257863 122846
rect 258022 122844 258028 122846
rect 258092 122844 258098 122908
rect 257797 122770 257863 122773
rect 258022 122770 258028 122772
rect 257797 122768 258028 122770
rect 257797 122712 257802 122768
rect 257858 122712 258028 122768
rect 257797 122710 258028 122712
rect 257797 122707 257863 122710
rect 258022 122708 258028 122710
rect 258092 122708 258098 122772
rect 256785 121818 256851 121821
rect 256785 121816 260084 121818
rect 256785 121760 256790 121816
rect 256846 121760 260084 121816
rect 256785 121758 260084 121760
rect 256785 121755 256851 121758
rect 345422 121138 345428 121140
rect 343804 121078 345428 121138
rect 345422 121076 345428 121078
rect 345492 121076 345498 121140
rect 260054 116106 260114 117028
rect 345013 116378 345079 116381
rect 343804 116376 345079 116378
rect 343804 116320 345018 116376
rect 345074 116320 345079 116376
rect 343804 116318 345079 116320
rect 345013 116315 345079 116318
rect 238710 116046 260114 116106
rect 237046 115908 237052 115972
rect 237116 115970 237122 115972
rect 238710 115970 238770 116046
rect 237116 115910 238770 115970
rect 237116 115908 237122 115910
rect 257797 113250 257863 113253
rect 258022 113250 258028 113252
rect 257797 113248 258028 113250
rect 257797 113192 257802 113248
rect 257858 113192 258028 113248
rect 257797 113190 258028 113192
rect 257797 113187 257863 113190
rect 258022 113188 258028 113190
rect 258092 113188 258098 113252
rect 257797 113114 257863 113117
rect 258022 113114 258028 113116
rect 257797 113112 258028 113114
rect 257797 113056 257802 113112
rect 257858 113056 258028 113112
rect 257797 113054 258028 113056
rect 257797 113051 257863 113054
rect 258022 113052 258028 113054
rect 258092 113052 258098 113116
rect 256785 112978 256851 112981
rect 256785 112976 260084 112978
rect 256785 112920 256790 112976
rect 256846 112920 260084 112976
rect 256785 112918 260084 112920
rect 256785 112915 256851 112918
rect 580441 112842 580507 112845
rect 583520 112842 584960 112932
rect 580441 112840 584960 112842
rect 580441 112784 580446 112840
rect 580502 112784 584960 112840
rect 580441 112782 584960 112784
rect 580441 112779 580507 112782
rect 583520 112692 584960 112782
rect 345381 112298 345447 112301
rect 343804 112296 345447 112298
rect 343804 112240 345386 112296
rect 345442 112240 345447 112296
rect 343804 112238 345447 112240
rect 345381 112235 345447 112238
rect -960 110666 480 110756
rect 3601 110666 3667 110669
rect -960 110664 3667 110666
rect -960 110608 3606 110664
rect 3662 110608 3667 110664
rect -960 110606 3667 110608
rect -960 110516 480 110606
rect 3601 110603 3667 110606
rect 238518 107612 238524 107676
rect 238588 107674 238594 107676
rect 260054 107674 260114 108188
rect 238588 107614 260114 107674
rect 238588 107612 238594 107614
rect 345197 107538 345263 107541
rect 343804 107536 345263 107538
rect 343804 107480 345202 107536
rect 345258 107480 345263 107536
rect 343804 107478 345263 107480
rect 345197 107475 345263 107478
rect 256785 104138 256851 104141
rect 256785 104136 260084 104138
rect 256785 104080 256790 104136
rect 256846 104080 260084 104136
rect 256785 104078 260084 104080
rect 256785 104075 256851 104078
rect 257797 103594 257863 103597
rect 258022 103594 258028 103596
rect 257797 103592 258028 103594
rect 257797 103536 257802 103592
rect 257858 103536 258028 103592
rect 257797 103534 258028 103536
rect 257797 103531 257863 103534
rect 258022 103532 258028 103534
rect 258092 103532 258098 103596
rect 257797 103458 257863 103461
rect 258022 103458 258028 103460
rect 257797 103456 258028 103458
rect 257797 103400 257802 103456
rect 257858 103400 258028 103456
rect 257797 103398 258028 103400
rect 257797 103395 257863 103398
rect 258022 103396 258028 103398
rect 258092 103396 258098 103460
rect 344093 103458 344159 103461
rect 343804 103456 344159 103458
rect 343804 103400 344098 103456
rect 344154 103400 344159 103456
rect 343804 103398 344159 103400
rect 344093 103395 344159 103398
rect 342294 100676 342300 100740
rect 342364 100738 342370 100740
rect 342805 100738 342871 100741
rect 342364 100736 342871 100738
rect 342364 100680 342810 100736
rect 342866 100680 342871 100736
rect 342364 100678 342871 100680
rect 342364 100676 342370 100678
rect 342805 100675 342871 100678
rect 579613 99514 579679 99517
rect 583520 99514 584960 99604
rect 579613 99512 584960 99514
rect 579613 99456 579618 99512
rect 579674 99456 584960 99512
rect 579613 99454 584960 99456
rect 579613 99451 579679 99454
rect 583520 99364 584960 99454
rect 233734 97820 233740 97884
rect 233804 97882 233810 97884
rect 288985 97882 289051 97885
rect 233804 97880 289051 97882
rect 233804 97824 288990 97880
rect 289046 97824 289051 97880
rect 233804 97822 289051 97824
rect 233804 97820 233810 97822
rect 288985 97819 289051 97822
rect 330845 97882 330911 97885
rect 345054 97882 345060 97884
rect 330845 97880 345060 97882
rect 330845 97824 330850 97880
rect 330906 97824 345060 97880
rect 330845 97822 345060 97824
rect 330845 97819 330911 97822
rect 345054 97820 345060 97822
rect 345124 97820 345130 97884
rect -960 97610 480 97700
rect 238334 97684 238340 97748
rect 238404 97746 238410 97748
rect 272241 97746 272307 97749
rect 238404 97744 272307 97746
rect 238404 97688 272246 97744
rect 272302 97688 272307 97744
rect 238404 97686 272307 97688
rect 238404 97684 238410 97686
rect 272241 97683 272307 97686
rect -960 97550 674 97610
rect -960 97474 480 97550
rect 614 97474 674 97550
rect 237230 97548 237236 97612
rect 237300 97610 237306 97612
rect 260005 97610 260071 97613
rect 237300 97608 260071 97610
rect 237300 97552 260010 97608
rect 260066 97552 260071 97608
rect 237300 97550 260071 97552
rect 237300 97548 237306 97550
rect 260005 97547 260071 97550
rect -960 97460 674 97474
rect 246 97414 674 97460
rect 246 96930 306 97414
rect 246 96870 6930 96930
rect 6870 96658 6930 96870
rect 235206 96658 235212 96660
rect 6870 96598 235212 96658
rect 235206 96596 235212 96598
rect 235276 96596 235282 96660
rect 257797 93938 257863 93941
rect 258022 93938 258028 93940
rect 257797 93936 258028 93938
rect 257797 93880 257802 93936
rect 257858 93880 258028 93936
rect 257797 93878 258028 93880
rect 257797 93875 257863 93878
rect 258022 93876 258028 93878
rect 258092 93876 258098 93940
rect 257981 93802 258047 93805
rect 257936 93800 258090 93802
rect 257936 93744 257986 93800
rect 258042 93744 258090 93800
rect 257936 93742 258090 93744
rect 257981 93739 258090 93742
rect 258030 93668 258090 93739
rect 258022 93604 258028 93668
rect 258092 93604 258098 93668
rect 580533 86186 580599 86189
rect 583520 86186 584960 86276
rect 580533 86184 584960 86186
rect 580533 86128 580538 86184
rect 580594 86128 584960 86184
rect 580533 86126 584960 86128
rect 580533 86123 580599 86126
rect 583520 86036 584960 86126
rect -960 84690 480 84780
rect 3325 84690 3391 84693
rect -960 84688 3391 84690
rect -960 84632 3330 84688
rect 3386 84632 3391 84688
rect -960 84630 3391 84632
rect -960 84540 480 84630
rect 3325 84627 3391 84630
rect 257981 84284 258047 84285
rect 257981 84282 258028 84284
rect 257936 84280 258028 84282
rect 258092 84282 258098 84284
rect 257936 84224 257986 84280
rect 257936 84222 258028 84224
rect 257981 84220 258028 84222
rect 258092 84222 258174 84282
rect 258092 84220 258098 84222
rect 257981 84219 258047 84220
rect 257981 84148 258047 84149
rect 257981 84146 258028 84148
rect 257936 84144 258028 84146
rect 258092 84146 258098 84148
rect 257936 84088 257986 84144
rect 257936 84086 258028 84088
rect 257981 84084 258028 84086
rect 258092 84086 258174 84146
rect 258092 84084 258098 84086
rect 257981 84083 258047 84084
rect 80053 80746 80119 80749
rect 251766 80746 251772 80748
rect 80053 80744 251772 80746
rect 80053 80688 80058 80744
rect 80114 80688 251772 80744
rect 80053 80686 251772 80688
rect 80053 80683 80119 80686
rect 251766 80684 251772 80686
rect 251836 80684 251842 80748
rect 27613 79386 27679 79389
rect 247166 79386 247172 79388
rect 27613 79384 247172 79386
rect 27613 79328 27618 79384
rect 27674 79328 247172 79384
rect 27613 79326 247172 79328
rect 27613 79323 27679 79326
rect 247166 79324 247172 79326
rect 247236 79324 247242 79388
rect 258022 74700 258028 74764
rect 258092 74700 258098 74764
rect 258030 74629 258090 74700
rect 257981 74626 258090 74629
rect 257936 74624 258090 74626
rect 257936 74568 257986 74624
rect 258042 74568 258090 74624
rect 257936 74566 258090 74568
rect 257981 74563 258047 74566
rect 257981 74492 258047 74493
rect 257981 74490 258028 74492
rect 257936 74488 258028 74490
rect 258092 74490 258098 74492
rect 257936 74432 257986 74488
rect 257936 74430 258028 74432
rect 257981 74428 258028 74430
rect 258092 74430 258174 74490
rect 258092 74428 258098 74430
rect 257981 74427 258047 74428
rect 580349 72994 580415 72997
rect 583520 72994 584960 73084
rect 580349 72992 584960 72994
rect 580349 72936 580354 72992
rect 580410 72936 584960 72992
rect 580349 72934 584960 72936
rect 580349 72931 580415 72934
rect 583520 72844 584960 72934
rect -960 71634 480 71724
rect 3325 71634 3391 71637
rect -960 71632 3391 71634
rect -960 71576 3330 71632
rect 3386 71576 3391 71632
rect -960 71574 3391 71576
rect -960 71484 480 71574
rect 3325 71571 3391 71574
rect 258022 65044 258028 65108
rect 258092 65044 258098 65108
rect 258030 64973 258090 65044
rect 257981 64970 258090 64973
rect 257936 64968 258090 64970
rect 257936 64912 257986 64968
rect 258042 64912 258090 64968
rect 257936 64910 258090 64912
rect 257981 64907 258047 64910
rect 257981 64834 258047 64837
rect 257936 64832 258090 64834
rect 257936 64776 257986 64832
rect 258042 64776 258090 64832
rect 257936 64774 258090 64776
rect 257981 64771 258090 64774
rect 258030 64700 258090 64771
rect 258022 64636 258028 64700
rect 258092 64636 258098 64700
rect 580206 59604 580212 59668
rect 580276 59666 580282 59668
rect 583520 59666 584960 59756
rect 580276 59606 584960 59666
rect 580276 59604 580282 59606
rect 583520 59516 584960 59606
rect -960 58578 480 58668
rect 3325 58578 3391 58581
rect -960 58576 3391 58578
rect -960 58520 3330 58576
rect 3386 58520 3391 58576
rect -960 58518 3391 58520
rect -960 58428 480 58518
rect 3325 58515 3391 58518
rect 257981 55316 258047 55317
rect 257981 55314 258028 55316
rect 257936 55312 258028 55314
rect 258092 55314 258098 55316
rect 257936 55256 257986 55312
rect 257936 55254 258028 55256
rect 257981 55252 258028 55254
rect 258092 55254 258174 55314
rect 258092 55252 258098 55254
rect 257981 55251 258047 55252
rect 257981 55178 258047 55181
rect 257936 55176 258090 55178
rect 257936 55120 257986 55176
rect 258042 55120 258090 55176
rect 257936 55118 258090 55120
rect 257981 55115 258090 55118
rect 258030 55044 258090 55115
rect 258022 54980 258028 55044
rect 258092 54980 258098 55044
rect 580257 46338 580323 46341
rect 583520 46338 584960 46428
rect 580257 46336 584960 46338
rect 580257 46280 580262 46336
rect 580318 46280 584960 46336
rect 580257 46278 584960 46280
rect 580257 46275 580323 46278
rect 583520 46188 584960 46278
rect 257981 45660 258047 45661
rect 257981 45658 258028 45660
rect 257936 45656 258028 45658
rect 258092 45658 258098 45660
rect -960 45522 480 45612
rect 257936 45600 257986 45656
rect 257936 45598 258028 45600
rect 257981 45596 258028 45598
rect 258092 45598 258174 45658
rect 258092 45596 258098 45598
rect 257981 45595 258047 45596
rect 3509 45522 3575 45525
rect 257981 45522 258047 45525
rect -960 45520 3575 45522
rect -960 45464 3514 45520
rect 3570 45464 3575 45520
rect -960 45462 3575 45464
rect 257936 45520 258090 45522
rect 257936 45464 257986 45520
rect 258042 45464 258090 45520
rect 257936 45462 258090 45464
rect -960 45372 480 45462
rect 3509 45459 3575 45462
rect 257981 45459 258090 45462
rect 258030 45388 258090 45459
rect 258022 45324 258028 45388
rect 258092 45324 258098 45388
rect 114553 44842 114619 44845
rect 254710 44842 254716 44844
rect 114553 44840 254716 44842
rect 114553 44784 114558 44840
rect 114614 44784 254716 44840
rect 114553 44782 254716 44784
rect 114553 44779 114619 44782
rect 254710 44780 254716 44782
rect 254780 44780 254786 44844
rect 257981 36004 258047 36005
rect 257981 36002 258028 36004
rect 257936 36000 258028 36002
rect 258092 36002 258098 36004
rect 257936 35944 257986 36000
rect 257936 35942 258028 35944
rect 257981 35940 258028 35942
rect 258092 35942 258174 36002
rect 258092 35940 258098 35942
rect 257981 35939 258047 35940
rect 257981 35866 258047 35869
rect 257936 35864 258090 35866
rect 257936 35808 257986 35864
rect 258042 35808 258090 35864
rect 257936 35806 258090 35808
rect 257981 35803 258090 35806
rect 258030 35732 258090 35803
rect 258022 35668 258028 35732
rect 258092 35668 258098 35732
rect 583520 33146 584960 33236
rect 583342 33086 584960 33146
rect 583342 33010 583402 33086
rect 583520 33010 584960 33086
rect 583342 32996 584960 33010
rect 583342 32950 583586 32996
rect -960 32466 480 32556
rect 3509 32466 3575 32469
rect -960 32464 3575 32466
rect -960 32408 3514 32464
rect 3570 32408 3575 32464
rect -960 32406 3575 32408
rect -960 32316 480 32406
rect 3509 32403 3575 32406
rect 346894 31724 346900 31788
rect 346964 31786 346970 31788
rect 583526 31786 583586 32950
rect 346964 31726 583586 31786
rect 346964 31724 346970 31726
rect 257981 26348 258047 26349
rect 257981 26346 258028 26348
rect 257936 26344 258028 26346
rect 258092 26346 258098 26348
rect 257936 26288 257986 26344
rect 257936 26286 258028 26288
rect 257981 26284 258028 26286
rect 258092 26286 258174 26346
rect 258092 26284 258098 26286
rect 257981 26283 258047 26284
rect 257981 26212 258047 26213
rect 257981 26210 258028 26212
rect 257936 26208 258028 26210
rect 258092 26210 258098 26212
rect 257936 26152 257986 26208
rect 257936 26150 258028 26152
rect 257981 26148 258028 26150
rect 258092 26150 258174 26210
rect 258092 26148 258098 26150
rect 257981 26147 258047 26148
rect 579705 19818 579771 19821
rect 583520 19818 584960 19908
rect 579705 19816 584960 19818
rect 579705 19760 579710 19816
rect 579766 19760 584960 19816
rect 579705 19758 584960 19760
rect 579705 19755 579771 19758
rect 583520 19668 584960 19758
rect -960 19410 480 19500
rect 3509 19410 3575 19413
rect -960 19408 3575 19410
rect -960 19352 3514 19408
rect 3570 19352 3575 19408
rect -960 19350 3575 19352
rect -960 19260 480 19350
rect 3509 19347 3575 19350
rect 258022 16764 258028 16828
rect 258092 16764 258098 16828
rect 258030 16693 258090 16764
rect 257981 16690 258090 16693
rect 257936 16688 258090 16690
rect 257936 16632 257986 16688
rect 258042 16632 258090 16688
rect 257936 16630 258090 16632
rect 257981 16627 258047 16630
rect 257981 16554 258047 16557
rect 257936 16552 258090 16554
rect 257936 16496 257986 16552
rect 258042 16496 258090 16552
rect 257936 16494 258090 16496
rect 257981 16491 258090 16494
rect 258030 16420 258090 16491
rect 258022 16356 258028 16420
rect 258092 16356 258098 16420
rect 77385 14514 77451 14517
rect 251582 14514 251588 14516
rect 77385 14512 251588 14514
rect 77385 14456 77390 14512
rect 77446 14456 251588 14512
rect 77385 14454 251588 14456
rect 77385 14451 77451 14454
rect 251582 14452 251588 14454
rect 251652 14452 251658 14516
rect 111609 13698 111675 13701
rect 254526 13698 254532 13700
rect 111609 13696 254532 13698
rect 111609 13640 111614 13696
rect 111670 13640 254532 13696
rect 111609 13638 254532 13640
rect 111609 13635 111675 13638
rect 254526 13636 254532 13638
rect 254596 13636 254602 13700
rect 59353 13562 59419 13565
rect 250110 13562 250116 13564
rect 59353 13560 250116 13562
rect 59353 13504 59358 13560
rect 59414 13504 250116 13560
rect 59353 13502 250116 13504
rect 59353 13499 59419 13502
rect 250110 13500 250116 13502
rect 250180 13500 250186 13564
rect 44265 13426 44331 13429
rect 248822 13426 248828 13428
rect 44265 13424 248828 13426
rect 44265 13368 44270 13424
rect 44326 13368 248828 13424
rect 44265 13366 248828 13368
rect 44265 13363 44331 13366
rect 248822 13364 248828 13366
rect 248892 13364 248898 13428
rect 40217 13290 40283 13293
rect 248638 13290 248644 13292
rect 40217 13288 248644 13290
rect 40217 13232 40222 13288
rect 40278 13232 248644 13288
rect 40217 13230 248644 13232
rect 40217 13227 40283 13230
rect 248638 13228 248644 13230
rect 248708 13228 248714 13292
rect 22553 13154 22619 13157
rect 247350 13154 247356 13156
rect 22553 13152 247356 13154
rect 22553 13096 22558 13152
rect 22614 13096 247356 13152
rect 22553 13094 247356 13096
rect 22553 13091 22619 13094
rect 247350 13092 247356 13094
rect 247420 13092 247426 13156
rect 8753 13018 8819 13021
rect 245878 13018 245884 13020
rect 8753 13016 245884 13018
rect 8753 12960 8758 13016
rect 8814 12960 245884 13016
rect 8753 12958 245884 12960
rect 8753 12955 8819 12958
rect 245878 12956 245884 12958
rect 245948 12956 245954 13020
rect 79225 10434 79291 10437
rect 251214 10434 251220 10436
rect 79225 10432 251220 10434
rect 79225 10376 79230 10432
rect 79286 10376 251220 10432
rect 79225 10374 251220 10376
rect 79225 10371 79291 10374
rect 251214 10372 251220 10374
rect 251284 10372 251290 10436
rect 75913 10298 75979 10301
rect 251398 10298 251404 10300
rect 75913 10296 251404 10298
rect 75913 10240 75918 10296
rect 75974 10240 251404 10296
rect 75913 10238 251404 10240
rect 75913 10235 75979 10238
rect 251398 10236 251404 10238
rect 251468 10236 251474 10300
rect 131757 9618 131823 9621
rect 255446 9618 255452 9620
rect 131757 9616 255452 9618
rect 131757 9560 131762 9616
rect 131818 9560 255452 9616
rect 131757 9558 255452 9560
rect 131757 9555 131823 9558
rect 255446 9556 255452 9558
rect 255516 9556 255522 9620
rect 54937 9482 55003 9485
rect 248597 9482 248663 9485
rect 54937 9480 248663 9482
rect 54937 9424 54942 9480
rect 54998 9424 248602 9480
rect 248658 9424 248663 9480
rect 54937 9422 248663 9424
rect 54937 9419 55003 9422
rect 248597 9419 248663 9422
rect 39573 9346 39639 9349
rect 247861 9346 247927 9349
rect 39573 9344 247927 9346
rect 39573 9288 39578 9344
rect 39634 9288 247866 9344
rect 247922 9288 247927 9344
rect 39573 9286 247927 9288
rect 39573 9283 39639 9286
rect 247861 9283 247927 9286
rect 32397 9210 32463 9213
rect 247953 9210 248019 9213
rect 32397 9208 248019 9210
rect 32397 9152 32402 9208
rect 32458 9152 247958 9208
rect 248014 9152 248019 9208
rect 32397 9150 248019 9152
rect 32397 9147 32463 9150
rect 247953 9147 248019 9150
rect 21817 9074 21883 9077
rect 245745 9074 245811 9077
rect 21817 9072 245811 9074
rect 21817 9016 21822 9072
rect 21878 9016 245750 9072
rect 245806 9016 245811 9072
rect 21817 9014 245811 9016
rect 21817 9011 21883 9014
rect 245745 9011 245811 9014
rect 17033 8938 17099 8941
rect 245837 8938 245903 8941
rect 17033 8936 245903 8938
rect 17033 8880 17038 8936
rect 17094 8880 245842 8936
rect 245898 8880 245903 8936
rect 17033 8878 245903 8880
rect 17033 8875 17099 8878
rect 245837 8875 245903 8878
rect 167177 7714 167243 7717
rect 259126 7714 259132 7716
rect 167177 7712 259132 7714
rect 167177 7656 167182 7712
rect 167238 7656 259132 7712
rect 167177 7654 259132 7656
rect 167177 7651 167243 7654
rect 259126 7652 259132 7654
rect 259196 7652 259202 7716
rect 96245 7578 96311 7581
rect 252686 7578 252692 7580
rect 96245 7576 252692 7578
rect 96245 7520 96250 7576
rect 96306 7520 252692 7576
rect 96245 7518 252692 7520
rect 96245 7515 96311 7518
rect 252686 7516 252692 7518
rect 252756 7516 252762 7580
rect 257981 7036 258047 7037
rect 257981 7034 258028 7036
rect 257936 7032 258028 7034
rect 258092 7034 258098 7036
rect 257936 6976 257986 7032
rect 257936 6974 258028 6976
rect 257981 6972 258028 6974
rect 258092 6974 258174 7034
rect 258092 6972 258098 6974
rect 257981 6971 258047 6972
rect 182909 6898 182975 6901
rect 254485 6898 254551 6901
rect 182909 6896 254551 6898
rect 182909 6840 182914 6896
rect 182970 6840 254490 6896
rect 254546 6840 254551 6896
rect 182909 6838 254551 6840
rect 182909 6835 182975 6838
rect 254485 6835 254551 6838
rect 169569 6762 169635 6765
rect 258022 6762 258028 6764
rect 169569 6760 258028 6762
rect 169569 6704 169574 6760
rect 169630 6704 258028 6760
rect 169569 6702 258028 6704
rect 169569 6699 169635 6702
rect 258022 6700 258028 6702
rect 258092 6700 258098 6764
rect 144729 6626 144795 6629
rect 256141 6626 256207 6629
rect 144729 6624 256207 6626
rect -960 6490 480 6580
rect 144729 6568 144734 6624
rect 144790 6568 256146 6624
rect 256202 6568 256207 6624
rect 144729 6566 256207 6568
rect 144729 6563 144795 6566
rect 256141 6563 256207 6566
rect 580165 6626 580231 6629
rect 583520 6626 584960 6716
rect 580165 6624 584960 6626
rect 580165 6568 580170 6624
rect 580226 6568 584960 6624
rect 580165 6566 584960 6568
rect 580165 6563 580231 6566
rect 3417 6490 3483 6493
rect -960 6488 3483 6490
rect -960 6432 3422 6488
rect 3478 6432 3483 6488
rect -960 6430 3483 6432
rect -960 6340 480 6430
rect 3417 6427 3483 6430
rect 119889 6490 119955 6493
rect 254761 6490 254827 6493
rect 119889 6488 254827 6490
rect 119889 6432 119894 6488
rect 119950 6432 254766 6488
rect 254822 6432 254827 6488
rect 583520 6476 584960 6566
rect 119889 6430 254827 6432
rect 119889 6427 119955 6430
rect 254761 6427 254827 6430
rect 89161 6354 89227 6357
rect 251725 6354 251791 6357
rect 89161 6352 251791 6354
rect 89161 6296 89166 6352
rect 89222 6296 251730 6352
rect 251786 6296 251791 6352
rect 89161 6294 251791 6296
rect 89161 6291 89227 6294
rect 251725 6291 251791 6294
rect 71497 6218 71563 6221
rect 249885 6218 249951 6221
rect 71497 6216 249951 6218
rect 71497 6160 71502 6216
rect 71558 6160 249890 6216
rect 249946 6160 249951 6216
rect 71497 6158 249951 6160
rect 71497 6155 71563 6158
rect 249885 6155 249951 6158
rect 157793 5130 157859 5133
rect 256734 5130 256740 5132
rect 157793 5128 256740 5130
rect 157793 5072 157798 5128
rect 157854 5072 256740 5128
rect 157793 5070 256740 5072
rect 157793 5067 157859 5070
rect 256734 5068 256740 5070
rect 256804 5068 256810 5132
rect 95141 4994 95207 4997
rect 252502 4994 252508 4996
rect 95141 4992 252508 4994
rect 95141 4936 95146 4992
rect 95202 4936 252508 4992
rect 95141 4934 252508 4936
rect 95141 4931 95207 4934
rect 252502 4932 252508 4934
rect 252572 4932 252578 4996
rect 6453 4858 6519 4861
rect 245694 4858 245700 4860
rect 6453 4856 245700 4858
rect 6453 4800 6458 4856
rect 6514 4800 245700 4856
rect 6453 4798 245700 4800
rect 6453 4795 6519 4798
rect 245694 4796 245700 4798
rect 245764 4796 245770 4860
rect 344185 4042 344251 4045
rect 335310 4040 344251 4042
rect 335310 3984 344190 4040
rect 344246 3984 344251 4040
rect 335310 3982 344251 3984
rect 260414 3844 260420 3908
rect 260484 3906 260490 3908
rect 274817 3906 274883 3909
rect 260484 3904 274883 3906
rect 260484 3848 274822 3904
rect 274878 3848 274883 3904
rect 260484 3846 274883 3848
rect 260484 3844 260490 3846
rect 274817 3843 274883 3846
rect 260598 3708 260604 3772
rect 260668 3770 260674 3772
rect 306741 3770 306807 3773
rect 260668 3768 306807 3770
rect 260668 3712 306746 3768
rect 306802 3712 306807 3768
rect 260668 3710 306807 3712
rect 260668 3708 260674 3710
rect 306741 3707 306807 3710
rect 257838 3572 257844 3636
rect 257908 3634 257914 3636
rect 310237 3634 310303 3637
rect 257908 3632 310303 3634
rect 257908 3576 310242 3632
rect 310298 3576 310303 3632
rect 257908 3574 310303 3576
rect 257908 3572 257914 3574
rect 310237 3571 310303 3574
rect 136449 3498 136515 3501
rect 255262 3498 255268 3500
rect 136449 3496 255268 3498
rect 136449 3440 136454 3496
rect 136510 3440 255268 3496
rect 136449 3438 255268 3440
rect 136449 3435 136515 3438
rect 255262 3436 255268 3438
rect 255332 3436 255338 3500
rect 257654 3436 257660 3500
rect 257724 3498 257730 3500
rect 313825 3498 313891 3501
rect 257724 3496 313891 3498
rect 257724 3440 313830 3496
rect 313886 3440 313891 3496
rect 257724 3438 313891 3440
rect 257724 3436 257730 3438
rect 313825 3435 313891 3438
rect 24209 3362 24275 3365
rect 243486 3362 243492 3364
rect 24209 3360 243492 3362
rect 24209 3304 24214 3360
rect 24270 3304 243492 3360
rect 24209 3302 243492 3304
rect 24209 3299 24275 3302
rect 243486 3300 243492 3302
rect 243556 3300 243562 3364
rect 255221 3362 255287 3365
rect 317321 3362 317387 3365
rect 255221 3360 317387 3362
rect 255221 3304 255226 3360
rect 255282 3304 317326 3360
rect 317382 3304 317387 3360
rect 255221 3302 317387 3304
rect 255221 3299 255287 3302
rect 317321 3299 317387 3302
rect 335077 3362 335143 3365
rect 335310 3362 335370 3982
rect 344185 3979 344251 3982
rect 343357 3906 343423 3909
rect 343357 3904 345030 3906
rect 343357 3848 343362 3904
rect 343418 3848 345030 3904
rect 343357 3846 345030 3848
rect 343357 3843 343423 3846
rect 339861 3770 339927 3773
rect 344970 3770 345030 3846
rect 349705 3770 349771 3773
rect 339861 3768 344754 3770
rect 339861 3712 339866 3768
rect 339922 3712 344754 3768
rect 339861 3710 344754 3712
rect 344970 3768 349771 3770
rect 344970 3712 349710 3768
rect 349766 3712 349771 3768
rect 344970 3710 349771 3712
rect 339861 3707 339927 3710
rect 338665 3634 338731 3637
rect 344461 3634 344527 3637
rect 338665 3632 344527 3634
rect 338665 3576 338670 3632
rect 338726 3576 344466 3632
rect 344522 3576 344527 3632
rect 338665 3574 344527 3576
rect 338665 3571 338731 3574
rect 344461 3571 344527 3574
rect 343582 3436 343588 3500
rect 343652 3498 343658 3500
rect 344553 3498 344619 3501
rect 343652 3496 344619 3498
rect 343652 3440 344558 3496
rect 344614 3440 344619 3496
rect 343652 3438 344619 3440
rect 344694 3498 344754 3710
rect 349705 3707 349771 3710
rect 344829 3634 344895 3637
rect 349429 3634 349495 3637
rect 344829 3632 349495 3634
rect 344829 3576 344834 3632
rect 344890 3576 349434 3632
rect 349490 3576 349495 3632
rect 344829 3574 349495 3576
rect 344829 3571 344895 3574
rect 349429 3571 349495 3574
rect 345289 3498 345355 3501
rect 344694 3496 345355 3498
rect 344694 3440 345294 3496
rect 345350 3440 345355 3496
rect 344694 3438 345355 3440
rect 343652 3436 343658 3438
rect 344553 3435 344619 3438
rect 345289 3435 345355 3438
rect 335077 3360 335370 3362
rect 335077 3304 335082 3360
rect 335138 3304 335370 3360
rect 335077 3302 335370 3304
rect 342161 3362 342227 3365
rect 346485 3362 346551 3365
rect 467465 3362 467531 3365
rect 342161 3360 346551 3362
rect 342161 3304 342166 3360
rect 342222 3304 346490 3360
rect 346546 3304 346551 3360
rect 342161 3302 346551 3304
rect 335077 3299 335143 3302
rect 342161 3299 342227 3302
rect 346485 3299 346551 3302
rect 354630 3360 467531 3362
rect 354630 3304 467470 3360
rect 467526 3304 467531 3360
rect 354630 3302 467531 3304
rect 340965 3226 341031 3229
rect 344829 3226 344895 3229
rect 340965 3224 344895 3226
rect 340965 3168 340970 3224
rect 341026 3168 344834 3224
rect 344890 3168 344895 3224
rect 340965 3166 344895 3168
rect 340965 3163 341031 3166
rect 344829 3163 344895 3166
rect 344962 3164 344968 3228
rect 345032 3226 345038 3228
rect 354630 3226 354690 3302
rect 467465 3299 467531 3302
rect 345032 3166 354690 3226
rect 345032 3164 345038 3166
rect 336273 3090 336339 3093
rect 347129 3090 347195 3093
rect 336273 3088 347195 3090
rect 336273 3032 336278 3088
rect 336334 3032 347134 3088
rect 347190 3032 347195 3088
rect 336273 3030 347195 3032
rect 336273 3027 336339 3030
rect 347129 3027 347195 3030
<< via3 >>
rect 114324 498204 114388 498268
rect 118924 498204 118988 498268
rect 123340 498204 123404 498268
rect 150572 498204 150636 498268
rect 124812 498068 124876 498132
rect 125732 498068 125796 498132
rect 397684 498068 397748 498132
rect 425468 498068 425532 498132
rect 410380 497660 410444 497724
rect 120028 497388 120092 497452
rect 399892 497252 399956 497316
rect 403388 497252 403452 497316
rect 398972 497116 399036 497180
rect 405228 496980 405292 497044
rect 113036 496904 113100 496908
rect 113036 496848 113086 496904
rect 113086 496848 113100 496904
rect 113036 496844 113100 496848
rect 115428 496904 115492 496908
rect 115428 496848 115478 496904
rect 115478 496848 115492 496904
rect 115428 496844 115492 496848
rect 117636 496844 117700 496908
rect 121132 496844 121196 496908
rect 122420 496844 122484 496908
rect 125364 496844 125428 496908
rect 130516 496844 130580 496908
rect 135484 496844 135548 496908
rect 140636 496904 140700 496908
rect 140636 496848 140686 496904
rect 140686 496848 140700 496904
rect 140636 496844 140700 496848
rect 145604 496844 145668 496908
rect 155540 496844 155604 496908
rect 160508 496844 160572 496908
rect 392900 496844 392964 496908
rect 394188 496844 394252 496908
rect 395292 496844 395356 496908
rect 400996 496844 401060 496908
rect 402100 496844 402164 496908
rect 404676 496844 404740 496908
rect 405780 496904 405844 496908
rect 405780 496848 405794 496904
rect 405794 496848 405844 496904
rect 405780 496844 405844 496848
rect 415532 496844 415596 496908
rect 420132 496844 420196 496908
rect 430436 496844 430500 496908
rect 435404 496844 435468 496908
rect 440556 496844 440620 496908
rect 233740 393408 233804 393412
rect 233740 393352 233790 393408
rect 233790 393352 233804 393408
rect 233740 393348 233804 393352
rect 239628 385052 239692 385116
rect 293356 384780 293420 384844
rect 296300 384780 296364 384844
rect 295012 384644 295076 384708
rect 238524 384508 238588 384572
rect 290780 384372 290844 384436
rect 345060 384236 345124 384300
rect 238156 384100 238220 384164
rect 235212 383964 235276 384028
rect 291332 383692 291396 383756
rect 296852 383284 296916 383348
rect 290596 382876 290660 382940
rect 342300 382740 342364 382804
rect 342852 382604 342916 382668
rect 293172 382468 293236 382532
rect 296116 382332 296180 382396
rect 283972 382120 284036 382124
rect 283972 382064 283976 382120
rect 283976 382064 284032 382120
rect 284032 382064 284036 382120
rect 237236 381788 237300 381852
rect 258764 381788 258828 381852
rect 273852 381848 273916 381852
rect 273852 381792 273902 381848
rect 273902 381792 273916 381848
rect 273852 381788 273916 381792
rect 276060 381848 276124 381852
rect 276060 381792 276110 381848
rect 276110 381792 276124 381848
rect 276060 381788 276124 381792
rect 280292 381788 280356 381852
rect 282500 381848 282564 381852
rect 283972 382060 284036 382064
rect 290964 382060 291028 382124
rect 298140 382060 298204 382124
rect 288756 381924 288820 381988
rect 288940 381924 289004 381988
rect 291148 381924 291212 381988
rect 293908 381924 293972 381988
rect 295748 381984 295812 381988
rect 295748 381928 295762 381984
rect 295762 381928 295812 381984
rect 295748 381924 295812 381928
rect 296484 381924 296548 381988
rect 282500 381792 282514 381848
rect 282514 381792 282564 381848
rect 282500 381788 282564 381792
rect 345244 381788 345308 381852
rect 580212 381516 580276 381580
rect 239996 381440 240060 381444
rect 239996 381384 240010 381440
rect 240010 381384 240060 381440
rect 239996 381380 240060 381384
rect 242388 381380 242452 381444
rect 245516 381440 245580 381444
rect 245516 381384 245530 381440
rect 245530 381384 245580 381440
rect 245516 381380 245580 381384
rect 346900 381380 346964 381444
rect 258764 381108 258828 381172
rect 280292 381108 280356 381172
rect 291700 381108 291764 381172
rect 242388 380972 242452 381036
rect 237052 380564 237116 380628
rect 273852 380564 273916 380628
rect 283972 380564 284036 380628
rect 276060 380428 276124 380492
rect 282500 380428 282564 380492
rect 245516 380292 245580 380356
rect 239996 380156 240060 380220
rect 296116 374036 296180 374100
rect 296668 374036 296732 374100
rect 296116 373900 296180 373964
rect 296668 373900 296732 373964
rect 296116 364380 296180 364444
rect 296668 364380 296732 364444
rect 296116 364244 296180 364308
rect 296668 364244 296732 364308
rect 238340 363428 238404 363492
rect 238892 363428 238956 363492
rect 296116 354724 296180 354788
rect 296668 354724 296732 354788
rect 296116 354588 296180 354652
rect 296668 354588 296732 354652
rect 296116 345068 296180 345132
rect 296668 345068 296732 345132
rect 296116 344932 296180 344996
rect 296668 344932 296732 344996
rect 238892 339900 238956 339964
rect 239628 339900 239692 339964
rect 245884 338132 245948 338196
rect 254532 338132 254596 338196
rect 255636 338132 255700 338196
rect 255820 337996 255884 338060
rect 266492 337996 266556 338060
rect 245700 337860 245764 337924
rect 246252 337724 246316 337788
rect 247172 337860 247236 337924
rect 248276 337860 248340 337924
rect 247356 337724 247420 337788
rect 250116 337860 250180 337924
rect 250300 337452 250364 337516
rect 251404 337860 251468 337924
rect 251772 337860 251836 337924
rect 252876 337920 252940 337924
rect 252876 337864 252880 337920
rect 252880 337864 252936 337920
rect 252936 337864 252940 337920
rect 252876 337860 252940 337864
rect 254164 337898 254168 337924
rect 254168 337898 254224 337924
rect 254224 337898 254228 337924
rect 254164 337860 254228 337898
rect 252692 337588 252756 337652
rect 254716 337860 254780 337924
rect 255452 337724 255516 337788
rect 257108 337860 257172 337924
rect 259132 337860 259196 337924
rect 259684 337860 259748 337924
rect 259684 337724 259748 337788
rect 251588 337316 251652 337380
rect 261156 337860 261220 337924
rect 260788 337588 260852 337652
rect 262260 337860 262324 337924
rect 262444 337860 262508 337924
rect 264100 337860 264164 337924
rect 263732 337784 263796 337788
rect 263732 337728 263736 337784
rect 263736 337728 263792 337784
rect 263792 337728 263796 337784
rect 263732 337724 263796 337728
rect 270172 337860 270236 337924
rect 272380 337920 272444 337924
rect 272380 337864 272384 337920
rect 272384 337864 272440 337920
rect 272440 337864 272444 337920
rect 270356 337784 270420 337788
rect 270356 337728 270406 337784
rect 270406 337728 270420 337784
rect 270356 337724 270420 337728
rect 272380 337860 272444 337864
rect 274036 337860 274100 337924
rect 274956 337860 275020 337924
rect 275876 337860 275940 337924
rect 276060 337860 276124 337924
rect 265572 337452 265636 337516
rect 274404 337724 274468 337788
rect 278636 337860 278700 337924
rect 279740 337860 279804 337924
rect 280844 337898 280848 337924
rect 280848 337898 280904 337924
rect 280904 337898 280908 337924
rect 280844 337860 280908 337898
rect 274772 337452 274836 337516
rect 279556 337588 279620 337652
rect 281580 337724 281644 337788
rect 282316 337920 282380 337924
rect 282316 337864 282320 337920
rect 282320 337864 282376 337920
rect 282376 337864 282380 337920
rect 282316 337860 282380 337864
rect 282500 337724 282564 337788
rect 284708 337860 284772 337924
rect 286364 337860 286428 337924
rect 290780 337996 290844 338060
rect 285444 337724 285508 337788
rect 286732 337784 286796 337788
rect 286732 337728 286736 337784
rect 286736 337728 286792 337784
rect 286792 337728 286796 337784
rect 286732 337724 286796 337728
rect 288204 337860 288268 337924
rect 288388 337898 288392 337924
rect 288392 337898 288448 337924
rect 288448 337898 288452 337924
rect 288388 337860 288452 337898
rect 287836 337724 287900 337788
rect 289492 337860 289556 337924
rect 289308 337724 289372 337788
rect 288940 337316 289004 337380
rect 282684 336772 282748 336836
rect 283420 336832 283484 336836
rect 283420 336776 283470 336832
rect 283470 336776 283484 336832
rect 283420 336772 283484 336776
rect 285076 336772 285140 336836
rect 263916 336696 263980 336700
rect 263916 336640 263930 336696
rect 263930 336640 263980 336696
rect 263916 336636 263980 336640
rect 266308 336636 266372 336700
rect 280844 336696 280908 336700
rect 280844 336640 280894 336696
rect 280894 336640 280908 336696
rect 280844 336636 280908 336640
rect 258028 336500 258092 336564
rect 281580 336500 281644 336564
rect 285444 336364 285508 336428
rect 254164 336228 254228 336292
rect 262628 336228 262692 336292
rect 272380 336152 272444 336156
rect 272380 336096 272430 336152
rect 272430 336096 272444 336152
rect 272380 336092 272444 336096
rect 277164 336016 277228 336020
rect 277164 335960 277178 336016
rect 277178 335960 277228 336016
rect 277164 335956 277228 335960
rect 282316 335956 282380 336020
rect 254716 335820 254780 335884
rect 255268 335820 255332 335884
rect 259500 335820 259564 335884
rect 262444 335820 262508 335884
rect 283604 335820 283668 335884
rect 259868 335684 259932 335748
rect 268148 335684 268212 335748
rect 248276 335548 248340 335612
rect 265204 335608 265268 335612
rect 265204 335552 265254 335608
rect 265254 335552 265268 335608
rect 265204 335548 265268 335552
rect 268332 335548 268396 335612
rect 283788 335548 283852 335612
rect 284892 335548 284956 335612
rect 265020 335472 265084 335476
rect 265020 335416 265070 335472
rect 265070 335416 265084 335472
rect 265020 335412 265084 335416
rect 265388 335472 265452 335476
rect 265388 335416 265438 335472
rect 265438 335416 265452 335472
rect 265388 335412 265452 335416
rect 268516 335412 268580 335476
rect 269068 335412 269132 335476
rect 271644 335412 271708 335476
rect 283420 335472 283484 335476
rect 283420 335416 283470 335472
rect 283470 335416 283484 335472
rect 283420 335412 283484 335416
rect 283972 335472 284036 335476
rect 283972 335416 283986 335472
rect 283986 335416 284036 335472
rect 283972 335412 284036 335416
rect 284156 335472 284220 335476
rect 284156 335416 284170 335472
rect 284170 335416 284220 335472
rect 284156 335412 284220 335416
rect 243492 335276 243556 335340
rect 256924 335276 256988 335340
rect 260972 335336 261036 335340
rect 260972 335280 261022 335336
rect 261022 335280 261036 335336
rect 260972 335276 261036 335280
rect 274772 335276 274836 335340
rect 274956 335336 275020 335340
rect 274956 335280 275006 335336
rect 275006 335280 275020 335336
rect 274956 335276 275020 335280
rect 296116 335412 296180 335476
rect 296668 335412 296732 335476
rect 286916 335200 286980 335204
rect 286916 335144 286930 335200
rect 286930 335144 286980 335200
rect 286916 335140 286980 335144
rect 296668 335140 296732 335204
rect 289308 335004 289372 335068
rect 246068 334732 246132 334796
rect 252508 334732 252572 334796
rect 256740 334732 256804 334796
rect 254900 334460 254964 334524
rect 259500 334460 259564 334524
rect 291332 333916 291396 333980
rect 344508 333780 344572 333844
rect 248644 333236 248708 333300
rect 251220 333296 251284 333300
rect 251220 333240 251270 333296
rect 251270 333240 251284 333296
rect 251220 333236 251284 333240
rect 274220 333236 274284 333300
rect 278452 333296 278516 333300
rect 278452 333240 278502 333296
rect 278502 333240 278516 333296
rect 278452 333236 278516 333240
rect 248828 333100 248892 333164
rect 254716 332828 254780 332892
rect 298140 332148 298204 332212
rect 260788 331876 260852 331940
rect 288204 331876 288268 331940
rect 289124 331740 289188 331804
rect 263548 331196 263612 331260
rect 264100 331196 264164 331260
rect 263548 331120 263612 331124
rect 263548 331064 263562 331120
rect 263562 331064 263612 331120
rect 263548 331060 263612 331064
rect 257108 330516 257172 330580
rect 284156 330516 284220 330580
rect 255820 330380 255884 330444
rect 284708 330380 284772 330444
rect 263916 328204 263980 328268
rect 256924 328068 256988 328132
rect 254900 327932 254964 327996
rect 252876 327796 252940 327860
rect 246252 327660 246316 327724
rect 284892 327660 284956 327724
rect 259868 326572 259932 326636
rect 255636 326436 255700 326500
rect 246068 326300 246132 326364
rect 265572 326300 265636 326364
rect 296668 325816 296732 325820
rect 296668 325760 296682 325816
rect 296682 325760 296732 325816
rect 296668 325756 296732 325760
rect 296668 325484 296732 325548
rect 263548 321600 263612 321604
rect 263548 321544 263562 321600
rect 263562 321544 263612 321600
rect 263548 321540 263612 321544
rect 274036 320724 274100 320788
rect 296668 316160 296732 316164
rect 296668 316104 296682 316160
rect 296682 316104 296732 316160
rect 296668 316100 296732 316104
rect 296668 316024 296732 316028
rect 296668 315968 296682 316024
rect 296682 315968 296732 316024
rect 296668 315964 296732 315968
rect 296668 306580 296732 306644
rect 296668 306368 296732 306372
rect 296668 306312 296682 306368
rect 296682 306312 296732 306368
rect 296668 306308 296732 306312
rect 296668 296924 296732 296988
rect 296668 296516 296732 296580
rect 296668 287192 296732 287196
rect 296668 287136 296682 287192
rect 296682 287136 296732 287192
rect 296668 287132 296732 287136
rect 296668 286860 296732 286924
rect 296668 277536 296732 277540
rect 296668 277480 296682 277536
rect 296682 277480 296732 277536
rect 296668 277476 296732 277480
rect 296668 277204 296732 277268
rect 296668 267880 296732 267884
rect 296668 267824 296682 267880
rect 296682 267824 296732 267880
rect 296668 267820 296732 267824
rect 296668 267744 296732 267748
rect 296668 267688 296682 267744
rect 296682 267688 296732 267744
rect 296668 267684 296732 267688
rect 296668 248432 296732 248436
rect 296668 248376 296682 248432
rect 296682 248376 296732 248432
rect 296668 248372 296732 248376
rect 296668 248296 296732 248300
rect 296668 248240 296682 248296
rect 296682 248240 296732 248296
rect 296668 248236 296732 248240
rect 296668 238852 296732 238916
rect 296668 238444 296732 238508
rect 296668 229120 296732 229124
rect 296668 229064 296682 229120
rect 296682 229064 296732 229120
rect 296668 229060 296732 229064
rect 296668 228788 296732 228852
rect 296668 219464 296732 219468
rect 296668 219408 296682 219464
rect 296682 219408 296732 219464
rect 296668 219404 296732 219408
rect 296668 219328 296732 219332
rect 296668 219272 296682 219328
rect 296682 219272 296732 219328
rect 296668 219268 296732 219272
rect 238156 214508 238220 214572
rect 296668 209884 296732 209948
rect 296668 209672 296732 209676
rect 296668 209616 296682 209672
rect 296682 209616 296732 209672
rect 296668 209612 296732 209616
rect 296668 200228 296732 200292
rect 296668 200016 296732 200020
rect 296668 199960 296682 200016
rect 296682 199960 296732 200016
rect 296668 199956 296732 199960
rect 293908 194516 293972 194580
rect 296668 190572 296732 190636
rect 296668 190164 296732 190228
rect 279740 186900 279804 186964
rect 296668 180840 296732 180844
rect 296668 180784 296682 180840
rect 296682 180784 296732 180840
rect 296668 180780 296732 180784
rect 296668 180508 296732 180572
rect 293356 179964 293420 180028
rect 250300 177244 250364 177308
rect 288020 177244 288084 177308
rect 276060 175884 276124 175948
rect 274220 174660 274284 174724
rect 283788 174524 283852 174588
rect 283972 173436 284036 173500
rect 286180 173300 286244 173364
rect 289308 173164 289372 173228
rect 296668 171184 296732 171188
rect 296668 171128 296682 171184
rect 296682 171128 296732 171184
rect 296668 171124 296732 171128
rect 296668 171048 296732 171052
rect 296668 170992 296682 171048
rect 296682 170992 296732 171048
rect 296668 170988 296732 170992
rect 295012 170444 295076 170508
rect 282500 170308 282564 170372
rect 278452 166500 278516 166564
rect 278636 166364 278700 166428
rect 279556 166228 279620 166292
rect 274404 165004 274468 165068
rect 275876 164868 275940 164932
rect 296852 163372 296916 163436
rect 285076 162284 285140 162348
rect 286732 162148 286796 162212
rect 289492 162012 289556 162076
rect 296852 161468 296916 161532
rect 296116 161332 296180 161396
rect 296484 161332 296548 161396
rect 345428 161332 345492 161396
rect 290964 161196 291028 161260
rect 268516 161060 268580 161124
rect 343588 161060 343652 161124
rect 262628 160924 262692 160988
rect 282684 160788 282748 160852
rect 287836 160652 287900 160716
rect 277164 159564 277228 159628
rect 265204 159428 265268 159492
rect 286916 159428 286980 159492
rect 263732 159292 263796 159356
rect 296300 159292 296364 159356
rect 265388 158748 265452 158812
rect 265020 158612 265084 158676
rect 295748 158612 295812 158676
rect 296668 158612 296732 158676
rect 291148 158476 291212 158540
rect 293172 158476 293236 158540
rect 288756 158340 288820 158404
rect 290596 158340 290660 158404
rect 266492 158204 266556 158268
rect 271644 158204 271708 158268
rect 263548 158068 263612 158132
rect 270172 158068 270236 158132
rect 262260 157932 262324 157996
rect 291700 157796 291764 157860
rect 344692 157388 344756 157452
rect 260972 156572 261036 156636
rect 283604 156572 283668 156636
rect 268332 155892 268396 155956
rect 257844 155756 257908 155820
rect 260420 155620 260484 155684
rect 284156 155620 284220 155684
rect 296116 155620 296180 155684
rect 261156 155484 261220 155548
rect 270356 155484 270420 155548
rect 259684 155348 259748 155412
rect 260604 155348 260668 155412
rect 259500 155212 259564 155276
rect 284156 155212 284220 155276
rect 266308 155076 266372 155140
rect 257660 153852 257724 153916
rect 269068 153852 269132 153916
rect 268148 153716 268212 153780
rect 257476 151812 257540 151876
rect 258028 151812 258092 151876
rect 257476 151676 257540 151740
rect 258028 151676 258092 151740
rect 343404 148276 343468 148340
rect 345244 142836 345308 142900
rect 257476 142156 257540 142220
rect 258028 142156 258092 142220
rect 258028 141884 258092 141948
rect 258028 132500 258092 132564
rect 258028 132364 258092 132428
rect 344692 129780 344756 129844
rect 258028 122844 258092 122908
rect 258028 122708 258092 122772
rect 345428 121076 345492 121140
rect 237052 115908 237116 115972
rect 258028 113188 258092 113252
rect 258028 113052 258092 113116
rect 238524 107612 238588 107676
rect 258028 103532 258092 103596
rect 258028 103396 258092 103460
rect 342300 100676 342364 100740
rect 233740 97820 233804 97884
rect 345060 97820 345124 97884
rect 238340 97684 238404 97748
rect 237236 97548 237300 97612
rect 235212 96596 235276 96660
rect 258028 93876 258092 93940
rect 258028 93604 258092 93668
rect 258028 84280 258092 84284
rect 258028 84224 258042 84280
rect 258042 84224 258092 84280
rect 258028 84220 258092 84224
rect 258028 84144 258092 84148
rect 258028 84088 258042 84144
rect 258042 84088 258092 84144
rect 258028 84084 258092 84088
rect 251772 80684 251836 80748
rect 247172 79324 247236 79388
rect 258028 74700 258092 74764
rect 258028 74488 258092 74492
rect 258028 74432 258042 74488
rect 258042 74432 258092 74488
rect 258028 74428 258092 74432
rect 258028 65044 258092 65108
rect 258028 64636 258092 64700
rect 580212 59604 580276 59668
rect 258028 55312 258092 55316
rect 258028 55256 258042 55312
rect 258042 55256 258092 55312
rect 258028 55252 258092 55256
rect 258028 54980 258092 55044
rect 258028 45656 258092 45660
rect 258028 45600 258042 45656
rect 258042 45600 258092 45656
rect 258028 45596 258092 45600
rect 258028 45324 258092 45388
rect 254716 44780 254780 44844
rect 258028 36000 258092 36004
rect 258028 35944 258042 36000
rect 258042 35944 258092 36000
rect 258028 35940 258092 35944
rect 258028 35668 258092 35732
rect 346900 31724 346964 31788
rect 258028 26344 258092 26348
rect 258028 26288 258042 26344
rect 258042 26288 258092 26344
rect 258028 26284 258092 26288
rect 258028 26208 258092 26212
rect 258028 26152 258042 26208
rect 258042 26152 258092 26208
rect 258028 26148 258092 26152
rect 258028 16764 258092 16828
rect 258028 16356 258092 16420
rect 251588 14452 251652 14516
rect 254532 13636 254596 13700
rect 250116 13500 250180 13564
rect 248828 13364 248892 13428
rect 248644 13228 248708 13292
rect 247356 13092 247420 13156
rect 245884 12956 245948 13020
rect 251220 10372 251284 10436
rect 251404 10236 251468 10300
rect 255452 9556 255516 9620
rect 259132 7652 259196 7716
rect 252692 7516 252756 7580
rect 258028 7032 258092 7036
rect 258028 6976 258042 7032
rect 258042 6976 258092 7032
rect 258028 6972 258092 6976
rect 258028 6700 258092 6764
rect 256740 5068 256804 5132
rect 252508 4932 252572 4996
rect 245700 4796 245764 4860
rect 260420 3844 260484 3908
rect 260604 3708 260668 3772
rect 257844 3572 257908 3636
rect 255268 3436 255332 3500
rect 257660 3436 257724 3500
rect 243492 3300 243556 3364
rect 343588 3436 343652 3500
rect 344968 3164 345032 3228
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 682954 -8106 711002
rect -8726 682718 -8694 682954
rect -8458 682718 -8374 682954
rect -8138 682718 -8106 682954
rect -8726 682634 -8106 682718
rect -8726 682398 -8694 682634
rect -8458 682398 -8374 682634
rect -8138 682398 -8106 682634
rect -8726 646954 -8106 682398
rect -8726 646718 -8694 646954
rect -8458 646718 -8374 646954
rect -8138 646718 -8106 646954
rect -8726 646634 -8106 646718
rect -8726 646398 -8694 646634
rect -8458 646398 -8374 646634
rect -8138 646398 -8106 646634
rect -8726 610954 -8106 646398
rect -8726 610718 -8694 610954
rect -8458 610718 -8374 610954
rect -8138 610718 -8106 610954
rect -8726 610634 -8106 610718
rect -8726 610398 -8694 610634
rect -8458 610398 -8374 610634
rect -8138 610398 -8106 610634
rect -8726 574954 -8106 610398
rect -8726 574718 -8694 574954
rect -8458 574718 -8374 574954
rect -8138 574718 -8106 574954
rect -8726 574634 -8106 574718
rect -8726 574398 -8694 574634
rect -8458 574398 -8374 574634
rect -8138 574398 -8106 574634
rect -8726 538954 -8106 574398
rect -8726 538718 -8694 538954
rect -8458 538718 -8374 538954
rect -8138 538718 -8106 538954
rect -8726 538634 -8106 538718
rect -8726 538398 -8694 538634
rect -8458 538398 -8374 538634
rect -8138 538398 -8106 538634
rect -8726 502954 -8106 538398
rect -8726 502718 -8694 502954
rect -8458 502718 -8374 502954
rect -8138 502718 -8106 502954
rect -8726 502634 -8106 502718
rect -8726 502398 -8694 502634
rect -8458 502398 -8374 502634
rect -8138 502398 -8106 502634
rect -8726 466954 -8106 502398
rect -8726 466718 -8694 466954
rect -8458 466718 -8374 466954
rect -8138 466718 -8106 466954
rect -8726 466634 -8106 466718
rect -8726 466398 -8694 466634
rect -8458 466398 -8374 466634
rect -8138 466398 -8106 466634
rect -8726 430954 -8106 466398
rect -8726 430718 -8694 430954
rect -8458 430718 -8374 430954
rect -8138 430718 -8106 430954
rect -8726 430634 -8106 430718
rect -8726 430398 -8694 430634
rect -8458 430398 -8374 430634
rect -8138 430398 -8106 430634
rect -8726 394954 -8106 430398
rect -8726 394718 -8694 394954
rect -8458 394718 -8374 394954
rect -8138 394718 -8106 394954
rect -8726 394634 -8106 394718
rect -8726 394398 -8694 394634
rect -8458 394398 -8374 394634
rect -8138 394398 -8106 394634
rect -8726 358954 -8106 394398
rect -8726 358718 -8694 358954
rect -8458 358718 -8374 358954
rect -8138 358718 -8106 358954
rect -8726 358634 -8106 358718
rect -8726 358398 -8694 358634
rect -8458 358398 -8374 358634
rect -8138 358398 -8106 358634
rect -8726 322954 -8106 358398
rect -8726 322718 -8694 322954
rect -8458 322718 -8374 322954
rect -8138 322718 -8106 322954
rect -8726 322634 -8106 322718
rect -8726 322398 -8694 322634
rect -8458 322398 -8374 322634
rect -8138 322398 -8106 322634
rect -8726 286954 -8106 322398
rect -8726 286718 -8694 286954
rect -8458 286718 -8374 286954
rect -8138 286718 -8106 286954
rect -8726 286634 -8106 286718
rect -8726 286398 -8694 286634
rect -8458 286398 -8374 286634
rect -8138 286398 -8106 286634
rect -8726 250954 -8106 286398
rect -8726 250718 -8694 250954
rect -8458 250718 -8374 250954
rect -8138 250718 -8106 250954
rect -8726 250634 -8106 250718
rect -8726 250398 -8694 250634
rect -8458 250398 -8374 250634
rect -8138 250398 -8106 250634
rect -8726 214954 -8106 250398
rect -8726 214718 -8694 214954
rect -8458 214718 -8374 214954
rect -8138 214718 -8106 214954
rect -8726 214634 -8106 214718
rect -8726 214398 -8694 214634
rect -8458 214398 -8374 214634
rect -8138 214398 -8106 214634
rect -8726 178954 -8106 214398
rect -8726 178718 -8694 178954
rect -8458 178718 -8374 178954
rect -8138 178718 -8106 178954
rect -8726 178634 -8106 178718
rect -8726 178398 -8694 178634
rect -8458 178398 -8374 178634
rect -8138 178398 -8106 178634
rect -8726 142954 -8106 178398
rect -8726 142718 -8694 142954
rect -8458 142718 -8374 142954
rect -8138 142718 -8106 142954
rect -8726 142634 -8106 142718
rect -8726 142398 -8694 142634
rect -8458 142398 -8374 142634
rect -8138 142398 -8106 142634
rect -8726 106954 -8106 142398
rect -8726 106718 -8694 106954
rect -8458 106718 -8374 106954
rect -8138 106718 -8106 106954
rect -8726 106634 -8106 106718
rect -8726 106398 -8694 106634
rect -8458 106398 -8374 106634
rect -8138 106398 -8106 106634
rect -8726 70954 -8106 106398
rect -8726 70718 -8694 70954
rect -8458 70718 -8374 70954
rect -8138 70718 -8106 70954
rect -8726 70634 -8106 70718
rect -8726 70398 -8694 70634
rect -8458 70398 -8374 70634
rect -8138 70398 -8106 70634
rect -8726 34954 -8106 70398
rect -8726 34718 -8694 34954
rect -8458 34718 -8374 34954
rect -8138 34718 -8106 34954
rect -8726 34634 -8106 34718
rect -8726 34398 -8694 34634
rect -8458 34398 -8374 34634
rect -8138 34398 -8106 34634
rect -8726 -7066 -8106 34398
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 678454 -7146 710042
rect -7766 678218 -7734 678454
rect -7498 678218 -7414 678454
rect -7178 678218 -7146 678454
rect -7766 678134 -7146 678218
rect -7766 677898 -7734 678134
rect -7498 677898 -7414 678134
rect -7178 677898 -7146 678134
rect -7766 642454 -7146 677898
rect -7766 642218 -7734 642454
rect -7498 642218 -7414 642454
rect -7178 642218 -7146 642454
rect -7766 642134 -7146 642218
rect -7766 641898 -7734 642134
rect -7498 641898 -7414 642134
rect -7178 641898 -7146 642134
rect -7766 606454 -7146 641898
rect -7766 606218 -7734 606454
rect -7498 606218 -7414 606454
rect -7178 606218 -7146 606454
rect -7766 606134 -7146 606218
rect -7766 605898 -7734 606134
rect -7498 605898 -7414 606134
rect -7178 605898 -7146 606134
rect -7766 570454 -7146 605898
rect -7766 570218 -7734 570454
rect -7498 570218 -7414 570454
rect -7178 570218 -7146 570454
rect -7766 570134 -7146 570218
rect -7766 569898 -7734 570134
rect -7498 569898 -7414 570134
rect -7178 569898 -7146 570134
rect -7766 534454 -7146 569898
rect -7766 534218 -7734 534454
rect -7498 534218 -7414 534454
rect -7178 534218 -7146 534454
rect -7766 534134 -7146 534218
rect -7766 533898 -7734 534134
rect -7498 533898 -7414 534134
rect -7178 533898 -7146 534134
rect -7766 498454 -7146 533898
rect -7766 498218 -7734 498454
rect -7498 498218 -7414 498454
rect -7178 498218 -7146 498454
rect -7766 498134 -7146 498218
rect -7766 497898 -7734 498134
rect -7498 497898 -7414 498134
rect -7178 497898 -7146 498134
rect -7766 462454 -7146 497898
rect -7766 462218 -7734 462454
rect -7498 462218 -7414 462454
rect -7178 462218 -7146 462454
rect -7766 462134 -7146 462218
rect -7766 461898 -7734 462134
rect -7498 461898 -7414 462134
rect -7178 461898 -7146 462134
rect -7766 426454 -7146 461898
rect -7766 426218 -7734 426454
rect -7498 426218 -7414 426454
rect -7178 426218 -7146 426454
rect -7766 426134 -7146 426218
rect -7766 425898 -7734 426134
rect -7498 425898 -7414 426134
rect -7178 425898 -7146 426134
rect -7766 390454 -7146 425898
rect -7766 390218 -7734 390454
rect -7498 390218 -7414 390454
rect -7178 390218 -7146 390454
rect -7766 390134 -7146 390218
rect -7766 389898 -7734 390134
rect -7498 389898 -7414 390134
rect -7178 389898 -7146 390134
rect -7766 354454 -7146 389898
rect -7766 354218 -7734 354454
rect -7498 354218 -7414 354454
rect -7178 354218 -7146 354454
rect -7766 354134 -7146 354218
rect -7766 353898 -7734 354134
rect -7498 353898 -7414 354134
rect -7178 353898 -7146 354134
rect -7766 318454 -7146 353898
rect -7766 318218 -7734 318454
rect -7498 318218 -7414 318454
rect -7178 318218 -7146 318454
rect -7766 318134 -7146 318218
rect -7766 317898 -7734 318134
rect -7498 317898 -7414 318134
rect -7178 317898 -7146 318134
rect -7766 282454 -7146 317898
rect -7766 282218 -7734 282454
rect -7498 282218 -7414 282454
rect -7178 282218 -7146 282454
rect -7766 282134 -7146 282218
rect -7766 281898 -7734 282134
rect -7498 281898 -7414 282134
rect -7178 281898 -7146 282134
rect -7766 246454 -7146 281898
rect -7766 246218 -7734 246454
rect -7498 246218 -7414 246454
rect -7178 246218 -7146 246454
rect -7766 246134 -7146 246218
rect -7766 245898 -7734 246134
rect -7498 245898 -7414 246134
rect -7178 245898 -7146 246134
rect -7766 210454 -7146 245898
rect -7766 210218 -7734 210454
rect -7498 210218 -7414 210454
rect -7178 210218 -7146 210454
rect -7766 210134 -7146 210218
rect -7766 209898 -7734 210134
rect -7498 209898 -7414 210134
rect -7178 209898 -7146 210134
rect -7766 174454 -7146 209898
rect -7766 174218 -7734 174454
rect -7498 174218 -7414 174454
rect -7178 174218 -7146 174454
rect -7766 174134 -7146 174218
rect -7766 173898 -7734 174134
rect -7498 173898 -7414 174134
rect -7178 173898 -7146 174134
rect -7766 138454 -7146 173898
rect -7766 138218 -7734 138454
rect -7498 138218 -7414 138454
rect -7178 138218 -7146 138454
rect -7766 138134 -7146 138218
rect -7766 137898 -7734 138134
rect -7498 137898 -7414 138134
rect -7178 137898 -7146 138134
rect -7766 102454 -7146 137898
rect -7766 102218 -7734 102454
rect -7498 102218 -7414 102454
rect -7178 102218 -7146 102454
rect -7766 102134 -7146 102218
rect -7766 101898 -7734 102134
rect -7498 101898 -7414 102134
rect -7178 101898 -7146 102134
rect -7766 66454 -7146 101898
rect -7766 66218 -7734 66454
rect -7498 66218 -7414 66454
rect -7178 66218 -7146 66454
rect -7766 66134 -7146 66218
rect -7766 65898 -7734 66134
rect -7498 65898 -7414 66134
rect -7178 65898 -7146 66134
rect -7766 30454 -7146 65898
rect -7766 30218 -7734 30454
rect -7498 30218 -7414 30454
rect -7178 30218 -7146 30454
rect -7766 30134 -7146 30218
rect -7766 29898 -7734 30134
rect -7498 29898 -7414 30134
rect -7178 29898 -7146 30134
rect -7766 -6106 -7146 29898
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 673954 -6186 709082
rect -6806 673718 -6774 673954
rect -6538 673718 -6454 673954
rect -6218 673718 -6186 673954
rect -6806 673634 -6186 673718
rect -6806 673398 -6774 673634
rect -6538 673398 -6454 673634
rect -6218 673398 -6186 673634
rect -6806 637954 -6186 673398
rect -6806 637718 -6774 637954
rect -6538 637718 -6454 637954
rect -6218 637718 -6186 637954
rect -6806 637634 -6186 637718
rect -6806 637398 -6774 637634
rect -6538 637398 -6454 637634
rect -6218 637398 -6186 637634
rect -6806 601954 -6186 637398
rect -6806 601718 -6774 601954
rect -6538 601718 -6454 601954
rect -6218 601718 -6186 601954
rect -6806 601634 -6186 601718
rect -6806 601398 -6774 601634
rect -6538 601398 -6454 601634
rect -6218 601398 -6186 601634
rect -6806 565954 -6186 601398
rect -6806 565718 -6774 565954
rect -6538 565718 -6454 565954
rect -6218 565718 -6186 565954
rect -6806 565634 -6186 565718
rect -6806 565398 -6774 565634
rect -6538 565398 -6454 565634
rect -6218 565398 -6186 565634
rect -6806 529954 -6186 565398
rect -6806 529718 -6774 529954
rect -6538 529718 -6454 529954
rect -6218 529718 -6186 529954
rect -6806 529634 -6186 529718
rect -6806 529398 -6774 529634
rect -6538 529398 -6454 529634
rect -6218 529398 -6186 529634
rect -6806 493954 -6186 529398
rect -6806 493718 -6774 493954
rect -6538 493718 -6454 493954
rect -6218 493718 -6186 493954
rect -6806 493634 -6186 493718
rect -6806 493398 -6774 493634
rect -6538 493398 -6454 493634
rect -6218 493398 -6186 493634
rect -6806 457954 -6186 493398
rect -6806 457718 -6774 457954
rect -6538 457718 -6454 457954
rect -6218 457718 -6186 457954
rect -6806 457634 -6186 457718
rect -6806 457398 -6774 457634
rect -6538 457398 -6454 457634
rect -6218 457398 -6186 457634
rect -6806 421954 -6186 457398
rect -6806 421718 -6774 421954
rect -6538 421718 -6454 421954
rect -6218 421718 -6186 421954
rect -6806 421634 -6186 421718
rect -6806 421398 -6774 421634
rect -6538 421398 -6454 421634
rect -6218 421398 -6186 421634
rect -6806 385954 -6186 421398
rect -6806 385718 -6774 385954
rect -6538 385718 -6454 385954
rect -6218 385718 -6186 385954
rect -6806 385634 -6186 385718
rect -6806 385398 -6774 385634
rect -6538 385398 -6454 385634
rect -6218 385398 -6186 385634
rect -6806 349954 -6186 385398
rect -6806 349718 -6774 349954
rect -6538 349718 -6454 349954
rect -6218 349718 -6186 349954
rect -6806 349634 -6186 349718
rect -6806 349398 -6774 349634
rect -6538 349398 -6454 349634
rect -6218 349398 -6186 349634
rect -6806 313954 -6186 349398
rect -6806 313718 -6774 313954
rect -6538 313718 -6454 313954
rect -6218 313718 -6186 313954
rect -6806 313634 -6186 313718
rect -6806 313398 -6774 313634
rect -6538 313398 -6454 313634
rect -6218 313398 -6186 313634
rect -6806 277954 -6186 313398
rect -6806 277718 -6774 277954
rect -6538 277718 -6454 277954
rect -6218 277718 -6186 277954
rect -6806 277634 -6186 277718
rect -6806 277398 -6774 277634
rect -6538 277398 -6454 277634
rect -6218 277398 -6186 277634
rect -6806 241954 -6186 277398
rect -6806 241718 -6774 241954
rect -6538 241718 -6454 241954
rect -6218 241718 -6186 241954
rect -6806 241634 -6186 241718
rect -6806 241398 -6774 241634
rect -6538 241398 -6454 241634
rect -6218 241398 -6186 241634
rect -6806 205954 -6186 241398
rect -6806 205718 -6774 205954
rect -6538 205718 -6454 205954
rect -6218 205718 -6186 205954
rect -6806 205634 -6186 205718
rect -6806 205398 -6774 205634
rect -6538 205398 -6454 205634
rect -6218 205398 -6186 205634
rect -6806 169954 -6186 205398
rect -6806 169718 -6774 169954
rect -6538 169718 -6454 169954
rect -6218 169718 -6186 169954
rect -6806 169634 -6186 169718
rect -6806 169398 -6774 169634
rect -6538 169398 -6454 169634
rect -6218 169398 -6186 169634
rect -6806 133954 -6186 169398
rect -6806 133718 -6774 133954
rect -6538 133718 -6454 133954
rect -6218 133718 -6186 133954
rect -6806 133634 -6186 133718
rect -6806 133398 -6774 133634
rect -6538 133398 -6454 133634
rect -6218 133398 -6186 133634
rect -6806 97954 -6186 133398
rect -6806 97718 -6774 97954
rect -6538 97718 -6454 97954
rect -6218 97718 -6186 97954
rect -6806 97634 -6186 97718
rect -6806 97398 -6774 97634
rect -6538 97398 -6454 97634
rect -6218 97398 -6186 97634
rect -6806 61954 -6186 97398
rect -6806 61718 -6774 61954
rect -6538 61718 -6454 61954
rect -6218 61718 -6186 61954
rect -6806 61634 -6186 61718
rect -6806 61398 -6774 61634
rect -6538 61398 -6454 61634
rect -6218 61398 -6186 61634
rect -6806 25954 -6186 61398
rect -6806 25718 -6774 25954
rect -6538 25718 -6454 25954
rect -6218 25718 -6186 25954
rect -6806 25634 -6186 25718
rect -6806 25398 -6774 25634
rect -6538 25398 -6454 25634
rect -6218 25398 -6186 25634
rect -6806 -5146 -6186 25398
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 669454 -5226 708122
rect -5846 669218 -5814 669454
rect -5578 669218 -5494 669454
rect -5258 669218 -5226 669454
rect -5846 669134 -5226 669218
rect -5846 668898 -5814 669134
rect -5578 668898 -5494 669134
rect -5258 668898 -5226 669134
rect -5846 633454 -5226 668898
rect -5846 633218 -5814 633454
rect -5578 633218 -5494 633454
rect -5258 633218 -5226 633454
rect -5846 633134 -5226 633218
rect -5846 632898 -5814 633134
rect -5578 632898 -5494 633134
rect -5258 632898 -5226 633134
rect -5846 597454 -5226 632898
rect -5846 597218 -5814 597454
rect -5578 597218 -5494 597454
rect -5258 597218 -5226 597454
rect -5846 597134 -5226 597218
rect -5846 596898 -5814 597134
rect -5578 596898 -5494 597134
rect -5258 596898 -5226 597134
rect -5846 561454 -5226 596898
rect -5846 561218 -5814 561454
rect -5578 561218 -5494 561454
rect -5258 561218 -5226 561454
rect -5846 561134 -5226 561218
rect -5846 560898 -5814 561134
rect -5578 560898 -5494 561134
rect -5258 560898 -5226 561134
rect -5846 525454 -5226 560898
rect -5846 525218 -5814 525454
rect -5578 525218 -5494 525454
rect -5258 525218 -5226 525454
rect -5846 525134 -5226 525218
rect -5846 524898 -5814 525134
rect -5578 524898 -5494 525134
rect -5258 524898 -5226 525134
rect -5846 489454 -5226 524898
rect -5846 489218 -5814 489454
rect -5578 489218 -5494 489454
rect -5258 489218 -5226 489454
rect -5846 489134 -5226 489218
rect -5846 488898 -5814 489134
rect -5578 488898 -5494 489134
rect -5258 488898 -5226 489134
rect -5846 453454 -5226 488898
rect -5846 453218 -5814 453454
rect -5578 453218 -5494 453454
rect -5258 453218 -5226 453454
rect -5846 453134 -5226 453218
rect -5846 452898 -5814 453134
rect -5578 452898 -5494 453134
rect -5258 452898 -5226 453134
rect -5846 417454 -5226 452898
rect -5846 417218 -5814 417454
rect -5578 417218 -5494 417454
rect -5258 417218 -5226 417454
rect -5846 417134 -5226 417218
rect -5846 416898 -5814 417134
rect -5578 416898 -5494 417134
rect -5258 416898 -5226 417134
rect -5846 381454 -5226 416898
rect -5846 381218 -5814 381454
rect -5578 381218 -5494 381454
rect -5258 381218 -5226 381454
rect -5846 381134 -5226 381218
rect -5846 380898 -5814 381134
rect -5578 380898 -5494 381134
rect -5258 380898 -5226 381134
rect -5846 345454 -5226 380898
rect -5846 345218 -5814 345454
rect -5578 345218 -5494 345454
rect -5258 345218 -5226 345454
rect -5846 345134 -5226 345218
rect -5846 344898 -5814 345134
rect -5578 344898 -5494 345134
rect -5258 344898 -5226 345134
rect -5846 309454 -5226 344898
rect -5846 309218 -5814 309454
rect -5578 309218 -5494 309454
rect -5258 309218 -5226 309454
rect -5846 309134 -5226 309218
rect -5846 308898 -5814 309134
rect -5578 308898 -5494 309134
rect -5258 308898 -5226 309134
rect -5846 273454 -5226 308898
rect -5846 273218 -5814 273454
rect -5578 273218 -5494 273454
rect -5258 273218 -5226 273454
rect -5846 273134 -5226 273218
rect -5846 272898 -5814 273134
rect -5578 272898 -5494 273134
rect -5258 272898 -5226 273134
rect -5846 237454 -5226 272898
rect -5846 237218 -5814 237454
rect -5578 237218 -5494 237454
rect -5258 237218 -5226 237454
rect -5846 237134 -5226 237218
rect -5846 236898 -5814 237134
rect -5578 236898 -5494 237134
rect -5258 236898 -5226 237134
rect -5846 201454 -5226 236898
rect -5846 201218 -5814 201454
rect -5578 201218 -5494 201454
rect -5258 201218 -5226 201454
rect -5846 201134 -5226 201218
rect -5846 200898 -5814 201134
rect -5578 200898 -5494 201134
rect -5258 200898 -5226 201134
rect -5846 165454 -5226 200898
rect -5846 165218 -5814 165454
rect -5578 165218 -5494 165454
rect -5258 165218 -5226 165454
rect -5846 165134 -5226 165218
rect -5846 164898 -5814 165134
rect -5578 164898 -5494 165134
rect -5258 164898 -5226 165134
rect -5846 129454 -5226 164898
rect -5846 129218 -5814 129454
rect -5578 129218 -5494 129454
rect -5258 129218 -5226 129454
rect -5846 129134 -5226 129218
rect -5846 128898 -5814 129134
rect -5578 128898 -5494 129134
rect -5258 128898 -5226 129134
rect -5846 93454 -5226 128898
rect -5846 93218 -5814 93454
rect -5578 93218 -5494 93454
rect -5258 93218 -5226 93454
rect -5846 93134 -5226 93218
rect -5846 92898 -5814 93134
rect -5578 92898 -5494 93134
rect -5258 92898 -5226 93134
rect -5846 57454 -5226 92898
rect -5846 57218 -5814 57454
rect -5578 57218 -5494 57454
rect -5258 57218 -5226 57454
rect -5846 57134 -5226 57218
rect -5846 56898 -5814 57134
rect -5578 56898 -5494 57134
rect -5258 56898 -5226 57134
rect -5846 21454 -5226 56898
rect -5846 21218 -5814 21454
rect -5578 21218 -5494 21454
rect -5258 21218 -5226 21454
rect -5846 21134 -5226 21218
rect -5846 20898 -5814 21134
rect -5578 20898 -5494 21134
rect -5258 20898 -5226 21134
rect -5846 -4186 -5226 20898
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 700954 -4266 707162
rect -4886 700718 -4854 700954
rect -4618 700718 -4534 700954
rect -4298 700718 -4266 700954
rect -4886 700634 -4266 700718
rect -4886 700398 -4854 700634
rect -4618 700398 -4534 700634
rect -4298 700398 -4266 700634
rect -4886 664954 -4266 700398
rect -4886 664718 -4854 664954
rect -4618 664718 -4534 664954
rect -4298 664718 -4266 664954
rect -4886 664634 -4266 664718
rect -4886 664398 -4854 664634
rect -4618 664398 -4534 664634
rect -4298 664398 -4266 664634
rect -4886 628954 -4266 664398
rect -4886 628718 -4854 628954
rect -4618 628718 -4534 628954
rect -4298 628718 -4266 628954
rect -4886 628634 -4266 628718
rect -4886 628398 -4854 628634
rect -4618 628398 -4534 628634
rect -4298 628398 -4266 628634
rect -4886 592954 -4266 628398
rect -4886 592718 -4854 592954
rect -4618 592718 -4534 592954
rect -4298 592718 -4266 592954
rect -4886 592634 -4266 592718
rect -4886 592398 -4854 592634
rect -4618 592398 -4534 592634
rect -4298 592398 -4266 592634
rect -4886 556954 -4266 592398
rect -4886 556718 -4854 556954
rect -4618 556718 -4534 556954
rect -4298 556718 -4266 556954
rect -4886 556634 -4266 556718
rect -4886 556398 -4854 556634
rect -4618 556398 -4534 556634
rect -4298 556398 -4266 556634
rect -4886 520954 -4266 556398
rect -4886 520718 -4854 520954
rect -4618 520718 -4534 520954
rect -4298 520718 -4266 520954
rect -4886 520634 -4266 520718
rect -4886 520398 -4854 520634
rect -4618 520398 -4534 520634
rect -4298 520398 -4266 520634
rect -4886 484954 -4266 520398
rect -4886 484718 -4854 484954
rect -4618 484718 -4534 484954
rect -4298 484718 -4266 484954
rect -4886 484634 -4266 484718
rect -4886 484398 -4854 484634
rect -4618 484398 -4534 484634
rect -4298 484398 -4266 484634
rect -4886 448954 -4266 484398
rect -4886 448718 -4854 448954
rect -4618 448718 -4534 448954
rect -4298 448718 -4266 448954
rect -4886 448634 -4266 448718
rect -4886 448398 -4854 448634
rect -4618 448398 -4534 448634
rect -4298 448398 -4266 448634
rect -4886 412954 -4266 448398
rect -4886 412718 -4854 412954
rect -4618 412718 -4534 412954
rect -4298 412718 -4266 412954
rect -4886 412634 -4266 412718
rect -4886 412398 -4854 412634
rect -4618 412398 -4534 412634
rect -4298 412398 -4266 412634
rect -4886 376954 -4266 412398
rect -4886 376718 -4854 376954
rect -4618 376718 -4534 376954
rect -4298 376718 -4266 376954
rect -4886 376634 -4266 376718
rect -4886 376398 -4854 376634
rect -4618 376398 -4534 376634
rect -4298 376398 -4266 376634
rect -4886 340954 -4266 376398
rect -4886 340718 -4854 340954
rect -4618 340718 -4534 340954
rect -4298 340718 -4266 340954
rect -4886 340634 -4266 340718
rect -4886 340398 -4854 340634
rect -4618 340398 -4534 340634
rect -4298 340398 -4266 340634
rect -4886 304954 -4266 340398
rect -4886 304718 -4854 304954
rect -4618 304718 -4534 304954
rect -4298 304718 -4266 304954
rect -4886 304634 -4266 304718
rect -4886 304398 -4854 304634
rect -4618 304398 -4534 304634
rect -4298 304398 -4266 304634
rect -4886 268954 -4266 304398
rect -4886 268718 -4854 268954
rect -4618 268718 -4534 268954
rect -4298 268718 -4266 268954
rect -4886 268634 -4266 268718
rect -4886 268398 -4854 268634
rect -4618 268398 -4534 268634
rect -4298 268398 -4266 268634
rect -4886 232954 -4266 268398
rect -4886 232718 -4854 232954
rect -4618 232718 -4534 232954
rect -4298 232718 -4266 232954
rect -4886 232634 -4266 232718
rect -4886 232398 -4854 232634
rect -4618 232398 -4534 232634
rect -4298 232398 -4266 232634
rect -4886 196954 -4266 232398
rect -4886 196718 -4854 196954
rect -4618 196718 -4534 196954
rect -4298 196718 -4266 196954
rect -4886 196634 -4266 196718
rect -4886 196398 -4854 196634
rect -4618 196398 -4534 196634
rect -4298 196398 -4266 196634
rect -4886 160954 -4266 196398
rect -4886 160718 -4854 160954
rect -4618 160718 -4534 160954
rect -4298 160718 -4266 160954
rect -4886 160634 -4266 160718
rect -4886 160398 -4854 160634
rect -4618 160398 -4534 160634
rect -4298 160398 -4266 160634
rect -4886 124954 -4266 160398
rect -4886 124718 -4854 124954
rect -4618 124718 -4534 124954
rect -4298 124718 -4266 124954
rect -4886 124634 -4266 124718
rect -4886 124398 -4854 124634
rect -4618 124398 -4534 124634
rect -4298 124398 -4266 124634
rect -4886 88954 -4266 124398
rect -4886 88718 -4854 88954
rect -4618 88718 -4534 88954
rect -4298 88718 -4266 88954
rect -4886 88634 -4266 88718
rect -4886 88398 -4854 88634
rect -4618 88398 -4534 88634
rect -4298 88398 -4266 88634
rect -4886 52954 -4266 88398
rect -4886 52718 -4854 52954
rect -4618 52718 -4534 52954
rect -4298 52718 -4266 52954
rect -4886 52634 -4266 52718
rect -4886 52398 -4854 52634
rect -4618 52398 -4534 52634
rect -4298 52398 -4266 52634
rect -4886 16954 -4266 52398
rect -4886 16718 -4854 16954
rect -4618 16718 -4534 16954
rect -4298 16718 -4266 16954
rect -4886 16634 -4266 16718
rect -4886 16398 -4854 16634
rect -4618 16398 -4534 16634
rect -4298 16398 -4266 16634
rect -4886 -3226 -4266 16398
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 696454 -3306 706202
rect -3926 696218 -3894 696454
rect -3658 696218 -3574 696454
rect -3338 696218 -3306 696454
rect -3926 696134 -3306 696218
rect -3926 695898 -3894 696134
rect -3658 695898 -3574 696134
rect -3338 695898 -3306 696134
rect -3926 660454 -3306 695898
rect -3926 660218 -3894 660454
rect -3658 660218 -3574 660454
rect -3338 660218 -3306 660454
rect -3926 660134 -3306 660218
rect -3926 659898 -3894 660134
rect -3658 659898 -3574 660134
rect -3338 659898 -3306 660134
rect -3926 624454 -3306 659898
rect -3926 624218 -3894 624454
rect -3658 624218 -3574 624454
rect -3338 624218 -3306 624454
rect -3926 624134 -3306 624218
rect -3926 623898 -3894 624134
rect -3658 623898 -3574 624134
rect -3338 623898 -3306 624134
rect -3926 588454 -3306 623898
rect -3926 588218 -3894 588454
rect -3658 588218 -3574 588454
rect -3338 588218 -3306 588454
rect -3926 588134 -3306 588218
rect -3926 587898 -3894 588134
rect -3658 587898 -3574 588134
rect -3338 587898 -3306 588134
rect -3926 552454 -3306 587898
rect -3926 552218 -3894 552454
rect -3658 552218 -3574 552454
rect -3338 552218 -3306 552454
rect -3926 552134 -3306 552218
rect -3926 551898 -3894 552134
rect -3658 551898 -3574 552134
rect -3338 551898 -3306 552134
rect -3926 516454 -3306 551898
rect -3926 516218 -3894 516454
rect -3658 516218 -3574 516454
rect -3338 516218 -3306 516454
rect -3926 516134 -3306 516218
rect -3926 515898 -3894 516134
rect -3658 515898 -3574 516134
rect -3338 515898 -3306 516134
rect -3926 480454 -3306 515898
rect -3926 480218 -3894 480454
rect -3658 480218 -3574 480454
rect -3338 480218 -3306 480454
rect -3926 480134 -3306 480218
rect -3926 479898 -3894 480134
rect -3658 479898 -3574 480134
rect -3338 479898 -3306 480134
rect -3926 444454 -3306 479898
rect -3926 444218 -3894 444454
rect -3658 444218 -3574 444454
rect -3338 444218 -3306 444454
rect -3926 444134 -3306 444218
rect -3926 443898 -3894 444134
rect -3658 443898 -3574 444134
rect -3338 443898 -3306 444134
rect -3926 408454 -3306 443898
rect -3926 408218 -3894 408454
rect -3658 408218 -3574 408454
rect -3338 408218 -3306 408454
rect -3926 408134 -3306 408218
rect -3926 407898 -3894 408134
rect -3658 407898 -3574 408134
rect -3338 407898 -3306 408134
rect -3926 372454 -3306 407898
rect -3926 372218 -3894 372454
rect -3658 372218 -3574 372454
rect -3338 372218 -3306 372454
rect -3926 372134 -3306 372218
rect -3926 371898 -3894 372134
rect -3658 371898 -3574 372134
rect -3338 371898 -3306 372134
rect -3926 336454 -3306 371898
rect -3926 336218 -3894 336454
rect -3658 336218 -3574 336454
rect -3338 336218 -3306 336454
rect -3926 336134 -3306 336218
rect -3926 335898 -3894 336134
rect -3658 335898 -3574 336134
rect -3338 335898 -3306 336134
rect -3926 300454 -3306 335898
rect -3926 300218 -3894 300454
rect -3658 300218 -3574 300454
rect -3338 300218 -3306 300454
rect -3926 300134 -3306 300218
rect -3926 299898 -3894 300134
rect -3658 299898 -3574 300134
rect -3338 299898 -3306 300134
rect -3926 264454 -3306 299898
rect -3926 264218 -3894 264454
rect -3658 264218 -3574 264454
rect -3338 264218 -3306 264454
rect -3926 264134 -3306 264218
rect -3926 263898 -3894 264134
rect -3658 263898 -3574 264134
rect -3338 263898 -3306 264134
rect -3926 228454 -3306 263898
rect -3926 228218 -3894 228454
rect -3658 228218 -3574 228454
rect -3338 228218 -3306 228454
rect -3926 228134 -3306 228218
rect -3926 227898 -3894 228134
rect -3658 227898 -3574 228134
rect -3338 227898 -3306 228134
rect -3926 192454 -3306 227898
rect -3926 192218 -3894 192454
rect -3658 192218 -3574 192454
rect -3338 192218 -3306 192454
rect -3926 192134 -3306 192218
rect -3926 191898 -3894 192134
rect -3658 191898 -3574 192134
rect -3338 191898 -3306 192134
rect -3926 156454 -3306 191898
rect -3926 156218 -3894 156454
rect -3658 156218 -3574 156454
rect -3338 156218 -3306 156454
rect -3926 156134 -3306 156218
rect -3926 155898 -3894 156134
rect -3658 155898 -3574 156134
rect -3338 155898 -3306 156134
rect -3926 120454 -3306 155898
rect -3926 120218 -3894 120454
rect -3658 120218 -3574 120454
rect -3338 120218 -3306 120454
rect -3926 120134 -3306 120218
rect -3926 119898 -3894 120134
rect -3658 119898 -3574 120134
rect -3338 119898 -3306 120134
rect -3926 84454 -3306 119898
rect -3926 84218 -3894 84454
rect -3658 84218 -3574 84454
rect -3338 84218 -3306 84454
rect -3926 84134 -3306 84218
rect -3926 83898 -3894 84134
rect -3658 83898 -3574 84134
rect -3338 83898 -3306 84134
rect -3926 48454 -3306 83898
rect -3926 48218 -3894 48454
rect -3658 48218 -3574 48454
rect -3338 48218 -3306 48454
rect -3926 48134 -3306 48218
rect -3926 47898 -3894 48134
rect -3658 47898 -3574 48134
rect -3338 47898 -3306 48134
rect -3926 12454 -3306 47898
rect -3926 12218 -3894 12454
rect -3658 12218 -3574 12454
rect -3338 12218 -3306 12454
rect -3926 12134 -3306 12218
rect -3926 11898 -3894 12134
rect -3658 11898 -3574 12134
rect -3338 11898 -3306 12134
rect -3926 -2266 -3306 11898
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 691954 -2346 705242
rect -2966 691718 -2934 691954
rect -2698 691718 -2614 691954
rect -2378 691718 -2346 691954
rect -2966 691634 -2346 691718
rect -2966 691398 -2934 691634
rect -2698 691398 -2614 691634
rect -2378 691398 -2346 691634
rect -2966 655954 -2346 691398
rect -2966 655718 -2934 655954
rect -2698 655718 -2614 655954
rect -2378 655718 -2346 655954
rect -2966 655634 -2346 655718
rect -2966 655398 -2934 655634
rect -2698 655398 -2614 655634
rect -2378 655398 -2346 655634
rect -2966 619954 -2346 655398
rect -2966 619718 -2934 619954
rect -2698 619718 -2614 619954
rect -2378 619718 -2346 619954
rect -2966 619634 -2346 619718
rect -2966 619398 -2934 619634
rect -2698 619398 -2614 619634
rect -2378 619398 -2346 619634
rect -2966 583954 -2346 619398
rect -2966 583718 -2934 583954
rect -2698 583718 -2614 583954
rect -2378 583718 -2346 583954
rect -2966 583634 -2346 583718
rect -2966 583398 -2934 583634
rect -2698 583398 -2614 583634
rect -2378 583398 -2346 583634
rect -2966 547954 -2346 583398
rect -2966 547718 -2934 547954
rect -2698 547718 -2614 547954
rect -2378 547718 -2346 547954
rect -2966 547634 -2346 547718
rect -2966 547398 -2934 547634
rect -2698 547398 -2614 547634
rect -2378 547398 -2346 547634
rect -2966 511954 -2346 547398
rect -2966 511718 -2934 511954
rect -2698 511718 -2614 511954
rect -2378 511718 -2346 511954
rect -2966 511634 -2346 511718
rect -2966 511398 -2934 511634
rect -2698 511398 -2614 511634
rect -2378 511398 -2346 511634
rect -2966 475954 -2346 511398
rect -2966 475718 -2934 475954
rect -2698 475718 -2614 475954
rect -2378 475718 -2346 475954
rect -2966 475634 -2346 475718
rect -2966 475398 -2934 475634
rect -2698 475398 -2614 475634
rect -2378 475398 -2346 475634
rect -2966 439954 -2346 475398
rect -2966 439718 -2934 439954
rect -2698 439718 -2614 439954
rect -2378 439718 -2346 439954
rect -2966 439634 -2346 439718
rect -2966 439398 -2934 439634
rect -2698 439398 -2614 439634
rect -2378 439398 -2346 439634
rect -2966 403954 -2346 439398
rect -2966 403718 -2934 403954
rect -2698 403718 -2614 403954
rect -2378 403718 -2346 403954
rect -2966 403634 -2346 403718
rect -2966 403398 -2934 403634
rect -2698 403398 -2614 403634
rect -2378 403398 -2346 403634
rect -2966 367954 -2346 403398
rect -2966 367718 -2934 367954
rect -2698 367718 -2614 367954
rect -2378 367718 -2346 367954
rect -2966 367634 -2346 367718
rect -2966 367398 -2934 367634
rect -2698 367398 -2614 367634
rect -2378 367398 -2346 367634
rect -2966 331954 -2346 367398
rect -2966 331718 -2934 331954
rect -2698 331718 -2614 331954
rect -2378 331718 -2346 331954
rect -2966 331634 -2346 331718
rect -2966 331398 -2934 331634
rect -2698 331398 -2614 331634
rect -2378 331398 -2346 331634
rect -2966 295954 -2346 331398
rect -2966 295718 -2934 295954
rect -2698 295718 -2614 295954
rect -2378 295718 -2346 295954
rect -2966 295634 -2346 295718
rect -2966 295398 -2934 295634
rect -2698 295398 -2614 295634
rect -2378 295398 -2346 295634
rect -2966 259954 -2346 295398
rect -2966 259718 -2934 259954
rect -2698 259718 -2614 259954
rect -2378 259718 -2346 259954
rect -2966 259634 -2346 259718
rect -2966 259398 -2934 259634
rect -2698 259398 -2614 259634
rect -2378 259398 -2346 259634
rect -2966 223954 -2346 259398
rect -2966 223718 -2934 223954
rect -2698 223718 -2614 223954
rect -2378 223718 -2346 223954
rect -2966 223634 -2346 223718
rect -2966 223398 -2934 223634
rect -2698 223398 -2614 223634
rect -2378 223398 -2346 223634
rect -2966 187954 -2346 223398
rect -2966 187718 -2934 187954
rect -2698 187718 -2614 187954
rect -2378 187718 -2346 187954
rect -2966 187634 -2346 187718
rect -2966 187398 -2934 187634
rect -2698 187398 -2614 187634
rect -2378 187398 -2346 187634
rect -2966 151954 -2346 187398
rect -2966 151718 -2934 151954
rect -2698 151718 -2614 151954
rect -2378 151718 -2346 151954
rect -2966 151634 -2346 151718
rect -2966 151398 -2934 151634
rect -2698 151398 -2614 151634
rect -2378 151398 -2346 151634
rect -2966 115954 -2346 151398
rect -2966 115718 -2934 115954
rect -2698 115718 -2614 115954
rect -2378 115718 -2346 115954
rect -2966 115634 -2346 115718
rect -2966 115398 -2934 115634
rect -2698 115398 -2614 115634
rect -2378 115398 -2346 115634
rect -2966 79954 -2346 115398
rect -2966 79718 -2934 79954
rect -2698 79718 -2614 79954
rect -2378 79718 -2346 79954
rect -2966 79634 -2346 79718
rect -2966 79398 -2934 79634
rect -2698 79398 -2614 79634
rect -2378 79398 -2346 79634
rect -2966 43954 -2346 79398
rect -2966 43718 -2934 43954
rect -2698 43718 -2614 43954
rect -2378 43718 -2346 43954
rect -2966 43634 -2346 43718
rect -2966 43398 -2934 43634
rect -2698 43398 -2614 43634
rect -2378 43398 -2346 43634
rect -2966 7954 -2346 43398
rect -2966 7718 -2934 7954
rect -2698 7718 -2614 7954
rect -2378 7718 -2346 7954
rect -2966 7634 -2346 7718
rect -2966 7398 -2934 7634
rect -2698 7398 -2614 7634
rect -2378 7398 -2346 7634
rect -2966 -1306 -2346 7398
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 711590
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 1794 -7654 2414 -902
rect 6294 705798 6914 711590
rect 6294 705562 6326 705798
rect 6562 705562 6646 705798
rect 6882 705562 6914 705798
rect 6294 705478 6914 705562
rect 6294 705242 6326 705478
rect 6562 705242 6646 705478
rect 6882 705242 6914 705478
rect 6294 691954 6914 705242
rect 6294 691718 6326 691954
rect 6562 691718 6646 691954
rect 6882 691718 6914 691954
rect 6294 691634 6914 691718
rect 6294 691398 6326 691634
rect 6562 691398 6646 691634
rect 6882 691398 6914 691634
rect 6294 655954 6914 691398
rect 6294 655718 6326 655954
rect 6562 655718 6646 655954
rect 6882 655718 6914 655954
rect 6294 655634 6914 655718
rect 6294 655398 6326 655634
rect 6562 655398 6646 655634
rect 6882 655398 6914 655634
rect 6294 619954 6914 655398
rect 6294 619718 6326 619954
rect 6562 619718 6646 619954
rect 6882 619718 6914 619954
rect 6294 619634 6914 619718
rect 6294 619398 6326 619634
rect 6562 619398 6646 619634
rect 6882 619398 6914 619634
rect 6294 583954 6914 619398
rect 6294 583718 6326 583954
rect 6562 583718 6646 583954
rect 6882 583718 6914 583954
rect 6294 583634 6914 583718
rect 6294 583398 6326 583634
rect 6562 583398 6646 583634
rect 6882 583398 6914 583634
rect 6294 547954 6914 583398
rect 6294 547718 6326 547954
rect 6562 547718 6646 547954
rect 6882 547718 6914 547954
rect 6294 547634 6914 547718
rect 6294 547398 6326 547634
rect 6562 547398 6646 547634
rect 6882 547398 6914 547634
rect 6294 511954 6914 547398
rect 6294 511718 6326 511954
rect 6562 511718 6646 511954
rect 6882 511718 6914 511954
rect 6294 511634 6914 511718
rect 6294 511398 6326 511634
rect 6562 511398 6646 511634
rect 6882 511398 6914 511634
rect 6294 475954 6914 511398
rect 6294 475718 6326 475954
rect 6562 475718 6646 475954
rect 6882 475718 6914 475954
rect 6294 475634 6914 475718
rect 6294 475398 6326 475634
rect 6562 475398 6646 475634
rect 6882 475398 6914 475634
rect 6294 439954 6914 475398
rect 6294 439718 6326 439954
rect 6562 439718 6646 439954
rect 6882 439718 6914 439954
rect 6294 439634 6914 439718
rect 6294 439398 6326 439634
rect 6562 439398 6646 439634
rect 6882 439398 6914 439634
rect 6294 403954 6914 439398
rect 6294 403718 6326 403954
rect 6562 403718 6646 403954
rect 6882 403718 6914 403954
rect 6294 403634 6914 403718
rect 6294 403398 6326 403634
rect 6562 403398 6646 403634
rect 6882 403398 6914 403634
rect 6294 367954 6914 403398
rect 6294 367718 6326 367954
rect 6562 367718 6646 367954
rect 6882 367718 6914 367954
rect 6294 367634 6914 367718
rect 6294 367398 6326 367634
rect 6562 367398 6646 367634
rect 6882 367398 6914 367634
rect 6294 331954 6914 367398
rect 6294 331718 6326 331954
rect 6562 331718 6646 331954
rect 6882 331718 6914 331954
rect 6294 331634 6914 331718
rect 6294 331398 6326 331634
rect 6562 331398 6646 331634
rect 6882 331398 6914 331634
rect 6294 295954 6914 331398
rect 6294 295718 6326 295954
rect 6562 295718 6646 295954
rect 6882 295718 6914 295954
rect 6294 295634 6914 295718
rect 6294 295398 6326 295634
rect 6562 295398 6646 295634
rect 6882 295398 6914 295634
rect 6294 259954 6914 295398
rect 6294 259718 6326 259954
rect 6562 259718 6646 259954
rect 6882 259718 6914 259954
rect 6294 259634 6914 259718
rect 6294 259398 6326 259634
rect 6562 259398 6646 259634
rect 6882 259398 6914 259634
rect 6294 223954 6914 259398
rect 6294 223718 6326 223954
rect 6562 223718 6646 223954
rect 6882 223718 6914 223954
rect 6294 223634 6914 223718
rect 6294 223398 6326 223634
rect 6562 223398 6646 223634
rect 6882 223398 6914 223634
rect 6294 187954 6914 223398
rect 6294 187718 6326 187954
rect 6562 187718 6646 187954
rect 6882 187718 6914 187954
rect 6294 187634 6914 187718
rect 6294 187398 6326 187634
rect 6562 187398 6646 187634
rect 6882 187398 6914 187634
rect 6294 151954 6914 187398
rect 6294 151718 6326 151954
rect 6562 151718 6646 151954
rect 6882 151718 6914 151954
rect 6294 151634 6914 151718
rect 6294 151398 6326 151634
rect 6562 151398 6646 151634
rect 6882 151398 6914 151634
rect 6294 115954 6914 151398
rect 6294 115718 6326 115954
rect 6562 115718 6646 115954
rect 6882 115718 6914 115954
rect 6294 115634 6914 115718
rect 6294 115398 6326 115634
rect 6562 115398 6646 115634
rect 6882 115398 6914 115634
rect 6294 79954 6914 115398
rect 6294 79718 6326 79954
rect 6562 79718 6646 79954
rect 6882 79718 6914 79954
rect 6294 79634 6914 79718
rect 6294 79398 6326 79634
rect 6562 79398 6646 79634
rect 6882 79398 6914 79634
rect 6294 43954 6914 79398
rect 6294 43718 6326 43954
rect 6562 43718 6646 43954
rect 6882 43718 6914 43954
rect 6294 43634 6914 43718
rect 6294 43398 6326 43634
rect 6562 43398 6646 43634
rect 6882 43398 6914 43634
rect 6294 7954 6914 43398
rect 6294 7718 6326 7954
rect 6562 7718 6646 7954
rect 6882 7718 6914 7954
rect 6294 7634 6914 7718
rect 6294 7398 6326 7634
rect 6562 7398 6646 7634
rect 6882 7398 6914 7634
rect 6294 -1306 6914 7398
rect 6294 -1542 6326 -1306
rect 6562 -1542 6646 -1306
rect 6882 -1542 6914 -1306
rect 6294 -1626 6914 -1542
rect 6294 -1862 6326 -1626
rect 6562 -1862 6646 -1626
rect 6882 -1862 6914 -1626
rect 6294 -7654 6914 -1862
rect 10794 706758 11414 711590
rect 10794 706522 10826 706758
rect 11062 706522 11146 706758
rect 11382 706522 11414 706758
rect 10794 706438 11414 706522
rect 10794 706202 10826 706438
rect 11062 706202 11146 706438
rect 11382 706202 11414 706438
rect 10794 696454 11414 706202
rect 10794 696218 10826 696454
rect 11062 696218 11146 696454
rect 11382 696218 11414 696454
rect 10794 696134 11414 696218
rect 10794 695898 10826 696134
rect 11062 695898 11146 696134
rect 11382 695898 11414 696134
rect 10794 660454 11414 695898
rect 10794 660218 10826 660454
rect 11062 660218 11146 660454
rect 11382 660218 11414 660454
rect 10794 660134 11414 660218
rect 10794 659898 10826 660134
rect 11062 659898 11146 660134
rect 11382 659898 11414 660134
rect 10794 624454 11414 659898
rect 10794 624218 10826 624454
rect 11062 624218 11146 624454
rect 11382 624218 11414 624454
rect 10794 624134 11414 624218
rect 10794 623898 10826 624134
rect 11062 623898 11146 624134
rect 11382 623898 11414 624134
rect 10794 588454 11414 623898
rect 10794 588218 10826 588454
rect 11062 588218 11146 588454
rect 11382 588218 11414 588454
rect 10794 588134 11414 588218
rect 10794 587898 10826 588134
rect 11062 587898 11146 588134
rect 11382 587898 11414 588134
rect 10794 552454 11414 587898
rect 10794 552218 10826 552454
rect 11062 552218 11146 552454
rect 11382 552218 11414 552454
rect 10794 552134 11414 552218
rect 10794 551898 10826 552134
rect 11062 551898 11146 552134
rect 11382 551898 11414 552134
rect 10794 516454 11414 551898
rect 10794 516218 10826 516454
rect 11062 516218 11146 516454
rect 11382 516218 11414 516454
rect 10794 516134 11414 516218
rect 10794 515898 10826 516134
rect 11062 515898 11146 516134
rect 11382 515898 11414 516134
rect 10794 480454 11414 515898
rect 10794 480218 10826 480454
rect 11062 480218 11146 480454
rect 11382 480218 11414 480454
rect 10794 480134 11414 480218
rect 10794 479898 10826 480134
rect 11062 479898 11146 480134
rect 11382 479898 11414 480134
rect 10794 444454 11414 479898
rect 10794 444218 10826 444454
rect 11062 444218 11146 444454
rect 11382 444218 11414 444454
rect 10794 444134 11414 444218
rect 10794 443898 10826 444134
rect 11062 443898 11146 444134
rect 11382 443898 11414 444134
rect 10794 408454 11414 443898
rect 10794 408218 10826 408454
rect 11062 408218 11146 408454
rect 11382 408218 11414 408454
rect 10794 408134 11414 408218
rect 10794 407898 10826 408134
rect 11062 407898 11146 408134
rect 11382 407898 11414 408134
rect 10794 372454 11414 407898
rect 10794 372218 10826 372454
rect 11062 372218 11146 372454
rect 11382 372218 11414 372454
rect 10794 372134 11414 372218
rect 10794 371898 10826 372134
rect 11062 371898 11146 372134
rect 11382 371898 11414 372134
rect 10794 336454 11414 371898
rect 10794 336218 10826 336454
rect 11062 336218 11146 336454
rect 11382 336218 11414 336454
rect 10794 336134 11414 336218
rect 10794 335898 10826 336134
rect 11062 335898 11146 336134
rect 11382 335898 11414 336134
rect 10794 300454 11414 335898
rect 10794 300218 10826 300454
rect 11062 300218 11146 300454
rect 11382 300218 11414 300454
rect 10794 300134 11414 300218
rect 10794 299898 10826 300134
rect 11062 299898 11146 300134
rect 11382 299898 11414 300134
rect 10794 264454 11414 299898
rect 10794 264218 10826 264454
rect 11062 264218 11146 264454
rect 11382 264218 11414 264454
rect 10794 264134 11414 264218
rect 10794 263898 10826 264134
rect 11062 263898 11146 264134
rect 11382 263898 11414 264134
rect 10794 228454 11414 263898
rect 10794 228218 10826 228454
rect 11062 228218 11146 228454
rect 11382 228218 11414 228454
rect 10794 228134 11414 228218
rect 10794 227898 10826 228134
rect 11062 227898 11146 228134
rect 11382 227898 11414 228134
rect 10794 192454 11414 227898
rect 10794 192218 10826 192454
rect 11062 192218 11146 192454
rect 11382 192218 11414 192454
rect 10794 192134 11414 192218
rect 10794 191898 10826 192134
rect 11062 191898 11146 192134
rect 11382 191898 11414 192134
rect 10794 156454 11414 191898
rect 10794 156218 10826 156454
rect 11062 156218 11146 156454
rect 11382 156218 11414 156454
rect 10794 156134 11414 156218
rect 10794 155898 10826 156134
rect 11062 155898 11146 156134
rect 11382 155898 11414 156134
rect 10794 120454 11414 155898
rect 10794 120218 10826 120454
rect 11062 120218 11146 120454
rect 11382 120218 11414 120454
rect 10794 120134 11414 120218
rect 10794 119898 10826 120134
rect 11062 119898 11146 120134
rect 11382 119898 11414 120134
rect 10794 84454 11414 119898
rect 10794 84218 10826 84454
rect 11062 84218 11146 84454
rect 11382 84218 11414 84454
rect 10794 84134 11414 84218
rect 10794 83898 10826 84134
rect 11062 83898 11146 84134
rect 11382 83898 11414 84134
rect 10794 48454 11414 83898
rect 10794 48218 10826 48454
rect 11062 48218 11146 48454
rect 11382 48218 11414 48454
rect 10794 48134 11414 48218
rect 10794 47898 10826 48134
rect 11062 47898 11146 48134
rect 11382 47898 11414 48134
rect 10794 12454 11414 47898
rect 10794 12218 10826 12454
rect 11062 12218 11146 12454
rect 11382 12218 11414 12454
rect 10794 12134 11414 12218
rect 10794 11898 10826 12134
rect 11062 11898 11146 12134
rect 11382 11898 11414 12134
rect 10794 -2266 11414 11898
rect 10794 -2502 10826 -2266
rect 11062 -2502 11146 -2266
rect 11382 -2502 11414 -2266
rect 10794 -2586 11414 -2502
rect 10794 -2822 10826 -2586
rect 11062 -2822 11146 -2586
rect 11382 -2822 11414 -2586
rect 10794 -7654 11414 -2822
rect 15294 707718 15914 711590
rect 15294 707482 15326 707718
rect 15562 707482 15646 707718
rect 15882 707482 15914 707718
rect 15294 707398 15914 707482
rect 15294 707162 15326 707398
rect 15562 707162 15646 707398
rect 15882 707162 15914 707398
rect 15294 700954 15914 707162
rect 15294 700718 15326 700954
rect 15562 700718 15646 700954
rect 15882 700718 15914 700954
rect 15294 700634 15914 700718
rect 15294 700398 15326 700634
rect 15562 700398 15646 700634
rect 15882 700398 15914 700634
rect 15294 664954 15914 700398
rect 15294 664718 15326 664954
rect 15562 664718 15646 664954
rect 15882 664718 15914 664954
rect 15294 664634 15914 664718
rect 15294 664398 15326 664634
rect 15562 664398 15646 664634
rect 15882 664398 15914 664634
rect 15294 628954 15914 664398
rect 15294 628718 15326 628954
rect 15562 628718 15646 628954
rect 15882 628718 15914 628954
rect 15294 628634 15914 628718
rect 15294 628398 15326 628634
rect 15562 628398 15646 628634
rect 15882 628398 15914 628634
rect 15294 592954 15914 628398
rect 15294 592718 15326 592954
rect 15562 592718 15646 592954
rect 15882 592718 15914 592954
rect 15294 592634 15914 592718
rect 15294 592398 15326 592634
rect 15562 592398 15646 592634
rect 15882 592398 15914 592634
rect 15294 556954 15914 592398
rect 15294 556718 15326 556954
rect 15562 556718 15646 556954
rect 15882 556718 15914 556954
rect 15294 556634 15914 556718
rect 15294 556398 15326 556634
rect 15562 556398 15646 556634
rect 15882 556398 15914 556634
rect 15294 520954 15914 556398
rect 15294 520718 15326 520954
rect 15562 520718 15646 520954
rect 15882 520718 15914 520954
rect 15294 520634 15914 520718
rect 15294 520398 15326 520634
rect 15562 520398 15646 520634
rect 15882 520398 15914 520634
rect 15294 484954 15914 520398
rect 15294 484718 15326 484954
rect 15562 484718 15646 484954
rect 15882 484718 15914 484954
rect 15294 484634 15914 484718
rect 15294 484398 15326 484634
rect 15562 484398 15646 484634
rect 15882 484398 15914 484634
rect 15294 448954 15914 484398
rect 15294 448718 15326 448954
rect 15562 448718 15646 448954
rect 15882 448718 15914 448954
rect 15294 448634 15914 448718
rect 15294 448398 15326 448634
rect 15562 448398 15646 448634
rect 15882 448398 15914 448634
rect 15294 412954 15914 448398
rect 15294 412718 15326 412954
rect 15562 412718 15646 412954
rect 15882 412718 15914 412954
rect 15294 412634 15914 412718
rect 15294 412398 15326 412634
rect 15562 412398 15646 412634
rect 15882 412398 15914 412634
rect 15294 376954 15914 412398
rect 15294 376718 15326 376954
rect 15562 376718 15646 376954
rect 15882 376718 15914 376954
rect 15294 376634 15914 376718
rect 15294 376398 15326 376634
rect 15562 376398 15646 376634
rect 15882 376398 15914 376634
rect 15294 340954 15914 376398
rect 15294 340718 15326 340954
rect 15562 340718 15646 340954
rect 15882 340718 15914 340954
rect 15294 340634 15914 340718
rect 15294 340398 15326 340634
rect 15562 340398 15646 340634
rect 15882 340398 15914 340634
rect 15294 304954 15914 340398
rect 15294 304718 15326 304954
rect 15562 304718 15646 304954
rect 15882 304718 15914 304954
rect 15294 304634 15914 304718
rect 15294 304398 15326 304634
rect 15562 304398 15646 304634
rect 15882 304398 15914 304634
rect 15294 268954 15914 304398
rect 15294 268718 15326 268954
rect 15562 268718 15646 268954
rect 15882 268718 15914 268954
rect 15294 268634 15914 268718
rect 15294 268398 15326 268634
rect 15562 268398 15646 268634
rect 15882 268398 15914 268634
rect 15294 232954 15914 268398
rect 15294 232718 15326 232954
rect 15562 232718 15646 232954
rect 15882 232718 15914 232954
rect 15294 232634 15914 232718
rect 15294 232398 15326 232634
rect 15562 232398 15646 232634
rect 15882 232398 15914 232634
rect 15294 196954 15914 232398
rect 15294 196718 15326 196954
rect 15562 196718 15646 196954
rect 15882 196718 15914 196954
rect 15294 196634 15914 196718
rect 15294 196398 15326 196634
rect 15562 196398 15646 196634
rect 15882 196398 15914 196634
rect 15294 160954 15914 196398
rect 15294 160718 15326 160954
rect 15562 160718 15646 160954
rect 15882 160718 15914 160954
rect 15294 160634 15914 160718
rect 15294 160398 15326 160634
rect 15562 160398 15646 160634
rect 15882 160398 15914 160634
rect 15294 124954 15914 160398
rect 15294 124718 15326 124954
rect 15562 124718 15646 124954
rect 15882 124718 15914 124954
rect 15294 124634 15914 124718
rect 15294 124398 15326 124634
rect 15562 124398 15646 124634
rect 15882 124398 15914 124634
rect 15294 88954 15914 124398
rect 15294 88718 15326 88954
rect 15562 88718 15646 88954
rect 15882 88718 15914 88954
rect 15294 88634 15914 88718
rect 15294 88398 15326 88634
rect 15562 88398 15646 88634
rect 15882 88398 15914 88634
rect 15294 52954 15914 88398
rect 15294 52718 15326 52954
rect 15562 52718 15646 52954
rect 15882 52718 15914 52954
rect 15294 52634 15914 52718
rect 15294 52398 15326 52634
rect 15562 52398 15646 52634
rect 15882 52398 15914 52634
rect 15294 16954 15914 52398
rect 15294 16718 15326 16954
rect 15562 16718 15646 16954
rect 15882 16718 15914 16954
rect 15294 16634 15914 16718
rect 15294 16398 15326 16634
rect 15562 16398 15646 16634
rect 15882 16398 15914 16634
rect 15294 -3226 15914 16398
rect 15294 -3462 15326 -3226
rect 15562 -3462 15646 -3226
rect 15882 -3462 15914 -3226
rect 15294 -3546 15914 -3462
rect 15294 -3782 15326 -3546
rect 15562 -3782 15646 -3546
rect 15882 -3782 15914 -3546
rect 15294 -7654 15914 -3782
rect 19794 708678 20414 711590
rect 19794 708442 19826 708678
rect 20062 708442 20146 708678
rect 20382 708442 20414 708678
rect 19794 708358 20414 708442
rect 19794 708122 19826 708358
rect 20062 708122 20146 708358
rect 20382 708122 20414 708358
rect 19794 669454 20414 708122
rect 19794 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 20414 669454
rect 19794 669134 20414 669218
rect 19794 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 20414 669134
rect 19794 633454 20414 668898
rect 19794 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 20414 633454
rect 19794 633134 20414 633218
rect 19794 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 20414 633134
rect 19794 597454 20414 632898
rect 19794 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 20414 597454
rect 19794 597134 20414 597218
rect 19794 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 20414 597134
rect 19794 561454 20414 596898
rect 19794 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 20414 561454
rect 19794 561134 20414 561218
rect 19794 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 20414 561134
rect 19794 525454 20414 560898
rect 19794 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 20414 525454
rect 19794 525134 20414 525218
rect 19794 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 20414 525134
rect 19794 489454 20414 524898
rect 19794 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 20414 489454
rect 19794 489134 20414 489218
rect 19794 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 20414 489134
rect 19794 453454 20414 488898
rect 19794 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 20414 453454
rect 19794 453134 20414 453218
rect 19794 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 20414 453134
rect 19794 417454 20414 452898
rect 19794 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 20414 417454
rect 19794 417134 20414 417218
rect 19794 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 20414 417134
rect 19794 381454 20414 416898
rect 19794 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 20414 381454
rect 19794 381134 20414 381218
rect 19794 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 20414 381134
rect 19794 345454 20414 380898
rect 19794 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 20414 345454
rect 19794 345134 20414 345218
rect 19794 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 20414 345134
rect 19794 309454 20414 344898
rect 19794 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 20414 309454
rect 19794 309134 20414 309218
rect 19794 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 20414 309134
rect 19794 273454 20414 308898
rect 19794 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 20414 273454
rect 19794 273134 20414 273218
rect 19794 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 20414 273134
rect 19794 237454 20414 272898
rect 19794 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 20414 237454
rect 19794 237134 20414 237218
rect 19794 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 20414 237134
rect 19794 201454 20414 236898
rect 19794 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 20414 201454
rect 19794 201134 20414 201218
rect 19794 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 20414 201134
rect 19794 165454 20414 200898
rect 19794 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 20414 165454
rect 19794 165134 20414 165218
rect 19794 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 20414 165134
rect 19794 129454 20414 164898
rect 19794 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 20414 129454
rect 19794 129134 20414 129218
rect 19794 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 20414 129134
rect 19794 93454 20414 128898
rect 19794 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 20414 93454
rect 19794 93134 20414 93218
rect 19794 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 20414 93134
rect 19794 57454 20414 92898
rect 19794 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 20414 57454
rect 19794 57134 20414 57218
rect 19794 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 20414 57134
rect 19794 21454 20414 56898
rect 19794 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 20414 21454
rect 19794 21134 20414 21218
rect 19794 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 20414 21134
rect 19794 -4186 20414 20898
rect 19794 -4422 19826 -4186
rect 20062 -4422 20146 -4186
rect 20382 -4422 20414 -4186
rect 19794 -4506 20414 -4422
rect 19794 -4742 19826 -4506
rect 20062 -4742 20146 -4506
rect 20382 -4742 20414 -4506
rect 19794 -7654 20414 -4742
rect 24294 709638 24914 711590
rect 24294 709402 24326 709638
rect 24562 709402 24646 709638
rect 24882 709402 24914 709638
rect 24294 709318 24914 709402
rect 24294 709082 24326 709318
rect 24562 709082 24646 709318
rect 24882 709082 24914 709318
rect 24294 673954 24914 709082
rect 24294 673718 24326 673954
rect 24562 673718 24646 673954
rect 24882 673718 24914 673954
rect 24294 673634 24914 673718
rect 24294 673398 24326 673634
rect 24562 673398 24646 673634
rect 24882 673398 24914 673634
rect 24294 637954 24914 673398
rect 24294 637718 24326 637954
rect 24562 637718 24646 637954
rect 24882 637718 24914 637954
rect 24294 637634 24914 637718
rect 24294 637398 24326 637634
rect 24562 637398 24646 637634
rect 24882 637398 24914 637634
rect 24294 601954 24914 637398
rect 24294 601718 24326 601954
rect 24562 601718 24646 601954
rect 24882 601718 24914 601954
rect 24294 601634 24914 601718
rect 24294 601398 24326 601634
rect 24562 601398 24646 601634
rect 24882 601398 24914 601634
rect 24294 565954 24914 601398
rect 24294 565718 24326 565954
rect 24562 565718 24646 565954
rect 24882 565718 24914 565954
rect 24294 565634 24914 565718
rect 24294 565398 24326 565634
rect 24562 565398 24646 565634
rect 24882 565398 24914 565634
rect 24294 529954 24914 565398
rect 24294 529718 24326 529954
rect 24562 529718 24646 529954
rect 24882 529718 24914 529954
rect 24294 529634 24914 529718
rect 24294 529398 24326 529634
rect 24562 529398 24646 529634
rect 24882 529398 24914 529634
rect 24294 493954 24914 529398
rect 24294 493718 24326 493954
rect 24562 493718 24646 493954
rect 24882 493718 24914 493954
rect 24294 493634 24914 493718
rect 24294 493398 24326 493634
rect 24562 493398 24646 493634
rect 24882 493398 24914 493634
rect 24294 457954 24914 493398
rect 24294 457718 24326 457954
rect 24562 457718 24646 457954
rect 24882 457718 24914 457954
rect 24294 457634 24914 457718
rect 24294 457398 24326 457634
rect 24562 457398 24646 457634
rect 24882 457398 24914 457634
rect 24294 421954 24914 457398
rect 24294 421718 24326 421954
rect 24562 421718 24646 421954
rect 24882 421718 24914 421954
rect 24294 421634 24914 421718
rect 24294 421398 24326 421634
rect 24562 421398 24646 421634
rect 24882 421398 24914 421634
rect 24294 385954 24914 421398
rect 24294 385718 24326 385954
rect 24562 385718 24646 385954
rect 24882 385718 24914 385954
rect 24294 385634 24914 385718
rect 24294 385398 24326 385634
rect 24562 385398 24646 385634
rect 24882 385398 24914 385634
rect 24294 349954 24914 385398
rect 24294 349718 24326 349954
rect 24562 349718 24646 349954
rect 24882 349718 24914 349954
rect 24294 349634 24914 349718
rect 24294 349398 24326 349634
rect 24562 349398 24646 349634
rect 24882 349398 24914 349634
rect 24294 313954 24914 349398
rect 24294 313718 24326 313954
rect 24562 313718 24646 313954
rect 24882 313718 24914 313954
rect 24294 313634 24914 313718
rect 24294 313398 24326 313634
rect 24562 313398 24646 313634
rect 24882 313398 24914 313634
rect 24294 277954 24914 313398
rect 24294 277718 24326 277954
rect 24562 277718 24646 277954
rect 24882 277718 24914 277954
rect 24294 277634 24914 277718
rect 24294 277398 24326 277634
rect 24562 277398 24646 277634
rect 24882 277398 24914 277634
rect 24294 241954 24914 277398
rect 24294 241718 24326 241954
rect 24562 241718 24646 241954
rect 24882 241718 24914 241954
rect 24294 241634 24914 241718
rect 24294 241398 24326 241634
rect 24562 241398 24646 241634
rect 24882 241398 24914 241634
rect 24294 205954 24914 241398
rect 24294 205718 24326 205954
rect 24562 205718 24646 205954
rect 24882 205718 24914 205954
rect 24294 205634 24914 205718
rect 24294 205398 24326 205634
rect 24562 205398 24646 205634
rect 24882 205398 24914 205634
rect 24294 169954 24914 205398
rect 24294 169718 24326 169954
rect 24562 169718 24646 169954
rect 24882 169718 24914 169954
rect 24294 169634 24914 169718
rect 24294 169398 24326 169634
rect 24562 169398 24646 169634
rect 24882 169398 24914 169634
rect 24294 133954 24914 169398
rect 24294 133718 24326 133954
rect 24562 133718 24646 133954
rect 24882 133718 24914 133954
rect 24294 133634 24914 133718
rect 24294 133398 24326 133634
rect 24562 133398 24646 133634
rect 24882 133398 24914 133634
rect 24294 97954 24914 133398
rect 24294 97718 24326 97954
rect 24562 97718 24646 97954
rect 24882 97718 24914 97954
rect 24294 97634 24914 97718
rect 24294 97398 24326 97634
rect 24562 97398 24646 97634
rect 24882 97398 24914 97634
rect 24294 61954 24914 97398
rect 24294 61718 24326 61954
rect 24562 61718 24646 61954
rect 24882 61718 24914 61954
rect 24294 61634 24914 61718
rect 24294 61398 24326 61634
rect 24562 61398 24646 61634
rect 24882 61398 24914 61634
rect 24294 25954 24914 61398
rect 24294 25718 24326 25954
rect 24562 25718 24646 25954
rect 24882 25718 24914 25954
rect 24294 25634 24914 25718
rect 24294 25398 24326 25634
rect 24562 25398 24646 25634
rect 24882 25398 24914 25634
rect 24294 -5146 24914 25398
rect 24294 -5382 24326 -5146
rect 24562 -5382 24646 -5146
rect 24882 -5382 24914 -5146
rect 24294 -5466 24914 -5382
rect 24294 -5702 24326 -5466
rect 24562 -5702 24646 -5466
rect 24882 -5702 24914 -5466
rect 24294 -7654 24914 -5702
rect 28794 710598 29414 711590
rect 28794 710362 28826 710598
rect 29062 710362 29146 710598
rect 29382 710362 29414 710598
rect 28794 710278 29414 710362
rect 28794 710042 28826 710278
rect 29062 710042 29146 710278
rect 29382 710042 29414 710278
rect 28794 678454 29414 710042
rect 28794 678218 28826 678454
rect 29062 678218 29146 678454
rect 29382 678218 29414 678454
rect 28794 678134 29414 678218
rect 28794 677898 28826 678134
rect 29062 677898 29146 678134
rect 29382 677898 29414 678134
rect 28794 642454 29414 677898
rect 28794 642218 28826 642454
rect 29062 642218 29146 642454
rect 29382 642218 29414 642454
rect 28794 642134 29414 642218
rect 28794 641898 28826 642134
rect 29062 641898 29146 642134
rect 29382 641898 29414 642134
rect 28794 606454 29414 641898
rect 28794 606218 28826 606454
rect 29062 606218 29146 606454
rect 29382 606218 29414 606454
rect 28794 606134 29414 606218
rect 28794 605898 28826 606134
rect 29062 605898 29146 606134
rect 29382 605898 29414 606134
rect 28794 570454 29414 605898
rect 28794 570218 28826 570454
rect 29062 570218 29146 570454
rect 29382 570218 29414 570454
rect 28794 570134 29414 570218
rect 28794 569898 28826 570134
rect 29062 569898 29146 570134
rect 29382 569898 29414 570134
rect 28794 534454 29414 569898
rect 28794 534218 28826 534454
rect 29062 534218 29146 534454
rect 29382 534218 29414 534454
rect 28794 534134 29414 534218
rect 28794 533898 28826 534134
rect 29062 533898 29146 534134
rect 29382 533898 29414 534134
rect 28794 498454 29414 533898
rect 28794 498218 28826 498454
rect 29062 498218 29146 498454
rect 29382 498218 29414 498454
rect 28794 498134 29414 498218
rect 28794 497898 28826 498134
rect 29062 497898 29146 498134
rect 29382 497898 29414 498134
rect 28794 462454 29414 497898
rect 28794 462218 28826 462454
rect 29062 462218 29146 462454
rect 29382 462218 29414 462454
rect 28794 462134 29414 462218
rect 28794 461898 28826 462134
rect 29062 461898 29146 462134
rect 29382 461898 29414 462134
rect 28794 426454 29414 461898
rect 28794 426218 28826 426454
rect 29062 426218 29146 426454
rect 29382 426218 29414 426454
rect 28794 426134 29414 426218
rect 28794 425898 28826 426134
rect 29062 425898 29146 426134
rect 29382 425898 29414 426134
rect 28794 390454 29414 425898
rect 28794 390218 28826 390454
rect 29062 390218 29146 390454
rect 29382 390218 29414 390454
rect 28794 390134 29414 390218
rect 28794 389898 28826 390134
rect 29062 389898 29146 390134
rect 29382 389898 29414 390134
rect 28794 354454 29414 389898
rect 28794 354218 28826 354454
rect 29062 354218 29146 354454
rect 29382 354218 29414 354454
rect 28794 354134 29414 354218
rect 28794 353898 28826 354134
rect 29062 353898 29146 354134
rect 29382 353898 29414 354134
rect 28794 318454 29414 353898
rect 28794 318218 28826 318454
rect 29062 318218 29146 318454
rect 29382 318218 29414 318454
rect 28794 318134 29414 318218
rect 28794 317898 28826 318134
rect 29062 317898 29146 318134
rect 29382 317898 29414 318134
rect 28794 282454 29414 317898
rect 28794 282218 28826 282454
rect 29062 282218 29146 282454
rect 29382 282218 29414 282454
rect 28794 282134 29414 282218
rect 28794 281898 28826 282134
rect 29062 281898 29146 282134
rect 29382 281898 29414 282134
rect 28794 246454 29414 281898
rect 28794 246218 28826 246454
rect 29062 246218 29146 246454
rect 29382 246218 29414 246454
rect 28794 246134 29414 246218
rect 28794 245898 28826 246134
rect 29062 245898 29146 246134
rect 29382 245898 29414 246134
rect 28794 210454 29414 245898
rect 28794 210218 28826 210454
rect 29062 210218 29146 210454
rect 29382 210218 29414 210454
rect 28794 210134 29414 210218
rect 28794 209898 28826 210134
rect 29062 209898 29146 210134
rect 29382 209898 29414 210134
rect 28794 174454 29414 209898
rect 28794 174218 28826 174454
rect 29062 174218 29146 174454
rect 29382 174218 29414 174454
rect 28794 174134 29414 174218
rect 28794 173898 28826 174134
rect 29062 173898 29146 174134
rect 29382 173898 29414 174134
rect 28794 138454 29414 173898
rect 28794 138218 28826 138454
rect 29062 138218 29146 138454
rect 29382 138218 29414 138454
rect 28794 138134 29414 138218
rect 28794 137898 28826 138134
rect 29062 137898 29146 138134
rect 29382 137898 29414 138134
rect 28794 102454 29414 137898
rect 28794 102218 28826 102454
rect 29062 102218 29146 102454
rect 29382 102218 29414 102454
rect 28794 102134 29414 102218
rect 28794 101898 28826 102134
rect 29062 101898 29146 102134
rect 29382 101898 29414 102134
rect 28794 66454 29414 101898
rect 28794 66218 28826 66454
rect 29062 66218 29146 66454
rect 29382 66218 29414 66454
rect 28794 66134 29414 66218
rect 28794 65898 28826 66134
rect 29062 65898 29146 66134
rect 29382 65898 29414 66134
rect 28794 30454 29414 65898
rect 28794 30218 28826 30454
rect 29062 30218 29146 30454
rect 29382 30218 29414 30454
rect 28794 30134 29414 30218
rect 28794 29898 28826 30134
rect 29062 29898 29146 30134
rect 29382 29898 29414 30134
rect 28794 -6106 29414 29898
rect 28794 -6342 28826 -6106
rect 29062 -6342 29146 -6106
rect 29382 -6342 29414 -6106
rect 28794 -6426 29414 -6342
rect 28794 -6662 28826 -6426
rect 29062 -6662 29146 -6426
rect 29382 -6662 29414 -6426
rect 28794 -7654 29414 -6662
rect 33294 711558 33914 711590
rect 33294 711322 33326 711558
rect 33562 711322 33646 711558
rect 33882 711322 33914 711558
rect 33294 711238 33914 711322
rect 33294 711002 33326 711238
rect 33562 711002 33646 711238
rect 33882 711002 33914 711238
rect 33294 682954 33914 711002
rect 33294 682718 33326 682954
rect 33562 682718 33646 682954
rect 33882 682718 33914 682954
rect 33294 682634 33914 682718
rect 33294 682398 33326 682634
rect 33562 682398 33646 682634
rect 33882 682398 33914 682634
rect 33294 646954 33914 682398
rect 33294 646718 33326 646954
rect 33562 646718 33646 646954
rect 33882 646718 33914 646954
rect 33294 646634 33914 646718
rect 33294 646398 33326 646634
rect 33562 646398 33646 646634
rect 33882 646398 33914 646634
rect 33294 610954 33914 646398
rect 33294 610718 33326 610954
rect 33562 610718 33646 610954
rect 33882 610718 33914 610954
rect 33294 610634 33914 610718
rect 33294 610398 33326 610634
rect 33562 610398 33646 610634
rect 33882 610398 33914 610634
rect 33294 574954 33914 610398
rect 33294 574718 33326 574954
rect 33562 574718 33646 574954
rect 33882 574718 33914 574954
rect 33294 574634 33914 574718
rect 33294 574398 33326 574634
rect 33562 574398 33646 574634
rect 33882 574398 33914 574634
rect 33294 538954 33914 574398
rect 33294 538718 33326 538954
rect 33562 538718 33646 538954
rect 33882 538718 33914 538954
rect 33294 538634 33914 538718
rect 33294 538398 33326 538634
rect 33562 538398 33646 538634
rect 33882 538398 33914 538634
rect 33294 502954 33914 538398
rect 33294 502718 33326 502954
rect 33562 502718 33646 502954
rect 33882 502718 33914 502954
rect 33294 502634 33914 502718
rect 33294 502398 33326 502634
rect 33562 502398 33646 502634
rect 33882 502398 33914 502634
rect 33294 466954 33914 502398
rect 33294 466718 33326 466954
rect 33562 466718 33646 466954
rect 33882 466718 33914 466954
rect 33294 466634 33914 466718
rect 33294 466398 33326 466634
rect 33562 466398 33646 466634
rect 33882 466398 33914 466634
rect 33294 430954 33914 466398
rect 33294 430718 33326 430954
rect 33562 430718 33646 430954
rect 33882 430718 33914 430954
rect 33294 430634 33914 430718
rect 33294 430398 33326 430634
rect 33562 430398 33646 430634
rect 33882 430398 33914 430634
rect 33294 394954 33914 430398
rect 33294 394718 33326 394954
rect 33562 394718 33646 394954
rect 33882 394718 33914 394954
rect 33294 394634 33914 394718
rect 33294 394398 33326 394634
rect 33562 394398 33646 394634
rect 33882 394398 33914 394634
rect 33294 358954 33914 394398
rect 33294 358718 33326 358954
rect 33562 358718 33646 358954
rect 33882 358718 33914 358954
rect 33294 358634 33914 358718
rect 33294 358398 33326 358634
rect 33562 358398 33646 358634
rect 33882 358398 33914 358634
rect 33294 322954 33914 358398
rect 33294 322718 33326 322954
rect 33562 322718 33646 322954
rect 33882 322718 33914 322954
rect 33294 322634 33914 322718
rect 33294 322398 33326 322634
rect 33562 322398 33646 322634
rect 33882 322398 33914 322634
rect 33294 286954 33914 322398
rect 33294 286718 33326 286954
rect 33562 286718 33646 286954
rect 33882 286718 33914 286954
rect 33294 286634 33914 286718
rect 33294 286398 33326 286634
rect 33562 286398 33646 286634
rect 33882 286398 33914 286634
rect 33294 250954 33914 286398
rect 33294 250718 33326 250954
rect 33562 250718 33646 250954
rect 33882 250718 33914 250954
rect 33294 250634 33914 250718
rect 33294 250398 33326 250634
rect 33562 250398 33646 250634
rect 33882 250398 33914 250634
rect 33294 214954 33914 250398
rect 33294 214718 33326 214954
rect 33562 214718 33646 214954
rect 33882 214718 33914 214954
rect 33294 214634 33914 214718
rect 33294 214398 33326 214634
rect 33562 214398 33646 214634
rect 33882 214398 33914 214634
rect 33294 178954 33914 214398
rect 33294 178718 33326 178954
rect 33562 178718 33646 178954
rect 33882 178718 33914 178954
rect 33294 178634 33914 178718
rect 33294 178398 33326 178634
rect 33562 178398 33646 178634
rect 33882 178398 33914 178634
rect 33294 142954 33914 178398
rect 33294 142718 33326 142954
rect 33562 142718 33646 142954
rect 33882 142718 33914 142954
rect 33294 142634 33914 142718
rect 33294 142398 33326 142634
rect 33562 142398 33646 142634
rect 33882 142398 33914 142634
rect 33294 106954 33914 142398
rect 33294 106718 33326 106954
rect 33562 106718 33646 106954
rect 33882 106718 33914 106954
rect 33294 106634 33914 106718
rect 33294 106398 33326 106634
rect 33562 106398 33646 106634
rect 33882 106398 33914 106634
rect 33294 70954 33914 106398
rect 33294 70718 33326 70954
rect 33562 70718 33646 70954
rect 33882 70718 33914 70954
rect 33294 70634 33914 70718
rect 33294 70398 33326 70634
rect 33562 70398 33646 70634
rect 33882 70398 33914 70634
rect 33294 34954 33914 70398
rect 33294 34718 33326 34954
rect 33562 34718 33646 34954
rect 33882 34718 33914 34954
rect 33294 34634 33914 34718
rect 33294 34398 33326 34634
rect 33562 34398 33646 34634
rect 33882 34398 33914 34634
rect 33294 -7066 33914 34398
rect 33294 -7302 33326 -7066
rect 33562 -7302 33646 -7066
rect 33882 -7302 33914 -7066
rect 33294 -7386 33914 -7302
rect 33294 -7622 33326 -7386
rect 33562 -7622 33646 -7386
rect 33882 -7622 33914 -7386
rect 33294 -7654 33914 -7622
rect 37794 704838 38414 711590
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 651454 38414 686898
rect 37794 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 38414 651454
rect 37794 651134 38414 651218
rect 37794 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 38414 651134
rect 37794 615454 38414 650898
rect 37794 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 38414 615454
rect 37794 615134 38414 615218
rect 37794 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 38414 615134
rect 37794 579454 38414 614898
rect 37794 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 38414 579454
rect 37794 579134 38414 579218
rect 37794 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 38414 579134
rect 37794 543454 38414 578898
rect 37794 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 38414 543454
rect 37794 543134 38414 543218
rect 37794 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 38414 543134
rect 37794 507454 38414 542898
rect 37794 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 38414 507454
rect 37794 507134 38414 507218
rect 37794 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 38414 507134
rect 37794 471454 38414 506898
rect 37794 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 38414 471454
rect 37794 471134 38414 471218
rect 37794 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 38414 471134
rect 37794 435454 38414 470898
rect 37794 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 38414 435454
rect 37794 435134 38414 435218
rect 37794 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 38414 435134
rect 37794 399454 38414 434898
rect 37794 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 38414 399454
rect 37794 399134 38414 399218
rect 37794 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 38414 399134
rect 37794 363454 38414 398898
rect 37794 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 38414 363454
rect 37794 363134 38414 363218
rect 37794 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 38414 363134
rect 37794 327454 38414 362898
rect 37794 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 38414 327454
rect 37794 327134 38414 327218
rect 37794 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 38414 327134
rect 37794 291454 38414 326898
rect 37794 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 38414 291454
rect 37794 291134 38414 291218
rect 37794 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 38414 291134
rect 37794 255454 38414 290898
rect 37794 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 38414 255454
rect 37794 255134 38414 255218
rect 37794 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 38414 255134
rect 37794 219454 38414 254898
rect 37794 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 38414 219454
rect 37794 219134 38414 219218
rect 37794 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 38414 219134
rect 37794 183454 38414 218898
rect 37794 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 38414 183454
rect 37794 183134 38414 183218
rect 37794 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 38414 183134
rect 37794 147454 38414 182898
rect 37794 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 38414 147454
rect 37794 147134 38414 147218
rect 37794 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 38414 147134
rect 37794 111454 38414 146898
rect 37794 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 38414 111454
rect 37794 111134 38414 111218
rect 37794 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 38414 111134
rect 37794 75454 38414 110898
rect 37794 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 38414 75454
rect 37794 75134 38414 75218
rect 37794 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 38414 75134
rect 37794 39454 38414 74898
rect 37794 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 38414 39454
rect 37794 39134 38414 39218
rect 37794 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 38414 39134
rect 37794 3454 38414 38898
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -7654 38414 -902
rect 42294 705798 42914 711590
rect 42294 705562 42326 705798
rect 42562 705562 42646 705798
rect 42882 705562 42914 705798
rect 42294 705478 42914 705562
rect 42294 705242 42326 705478
rect 42562 705242 42646 705478
rect 42882 705242 42914 705478
rect 42294 691954 42914 705242
rect 42294 691718 42326 691954
rect 42562 691718 42646 691954
rect 42882 691718 42914 691954
rect 42294 691634 42914 691718
rect 42294 691398 42326 691634
rect 42562 691398 42646 691634
rect 42882 691398 42914 691634
rect 42294 655954 42914 691398
rect 42294 655718 42326 655954
rect 42562 655718 42646 655954
rect 42882 655718 42914 655954
rect 42294 655634 42914 655718
rect 42294 655398 42326 655634
rect 42562 655398 42646 655634
rect 42882 655398 42914 655634
rect 42294 619954 42914 655398
rect 42294 619718 42326 619954
rect 42562 619718 42646 619954
rect 42882 619718 42914 619954
rect 42294 619634 42914 619718
rect 42294 619398 42326 619634
rect 42562 619398 42646 619634
rect 42882 619398 42914 619634
rect 42294 583954 42914 619398
rect 42294 583718 42326 583954
rect 42562 583718 42646 583954
rect 42882 583718 42914 583954
rect 42294 583634 42914 583718
rect 42294 583398 42326 583634
rect 42562 583398 42646 583634
rect 42882 583398 42914 583634
rect 42294 547954 42914 583398
rect 42294 547718 42326 547954
rect 42562 547718 42646 547954
rect 42882 547718 42914 547954
rect 42294 547634 42914 547718
rect 42294 547398 42326 547634
rect 42562 547398 42646 547634
rect 42882 547398 42914 547634
rect 42294 511954 42914 547398
rect 42294 511718 42326 511954
rect 42562 511718 42646 511954
rect 42882 511718 42914 511954
rect 42294 511634 42914 511718
rect 42294 511398 42326 511634
rect 42562 511398 42646 511634
rect 42882 511398 42914 511634
rect 42294 475954 42914 511398
rect 42294 475718 42326 475954
rect 42562 475718 42646 475954
rect 42882 475718 42914 475954
rect 42294 475634 42914 475718
rect 42294 475398 42326 475634
rect 42562 475398 42646 475634
rect 42882 475398 42914 475634
rect 42294 439954 42914 475398
rect 42294 439718 42326 439954
rect 42562 439718 42646 439954
rect 42882 439718 42914 439954
rect 42294 439634 42914 439718
rect 42294 439398 42326 439634
rect 42562 439398 42646 439634
rect 42882 439398 42914 439634
rect 42294 403954 42914 439398
rect 42294 403718 42326 403954
rect 42562 403718 42646 403954
rect 42882 403718 42914 403954
rect 42294 403634 42914 403718
rect 42294 403398 42326 403634
rect 42562 403398 42646 403634
rect 42882 403398 42914 403634
rect 42294 367954 42914 403398
rect 42294 367718 42326 367954
rect 42562 367718 42646 367954
rect 42882 367718 42914 367954
rect 42294 367634 42914 367718
rect 42294 367398 42326 367634
rect 42562 367398 42646 367634
rect 42882 367398 42914 367634
rect 42294 331954 42914 367398
rect 42294 331718 42326 331954
rect 42562 331718 42646 331954
rect 42882 331718 42914 331954
rect 42294 331634 42914 331718
rect 42294 331398 42326 331634
rect 42562 331398 42646 331634
rect 42882 331398 42914 331634
rect 42294 295954 42914 331398
rect 42294 295718 42326 295954
rect 42562 295718 42646 295954
rect 42882 295718 42914 295954
rect 42294 295634 42914 295718
rect 42294 295398 42326 295634
rect 42562 295398 42646 295634
rect 42882 295398 42914 295634
rect 42294 259954 42914 295398
rect 42294 259718 42326 259954
rect 42562 259718 42646 259954
rect 42882 259718 42914 259954
rect 42294 259634 42914 259718
rect 42294 259398 42326 259634
rect 42562 259398 42646 259634
rect 42882 259398 42914 259634
rect 42294 223954 42914 259398
rect 42294 223718 42326 223954
rect 42562 223718 42646 223954
rect 42882 223718 42914 223954
rect 42294 223634 42914 223718
rect 42294 223398 42326 223634
rect 42562 223398 42646 223634
rect 42882 223398 42914 223634
rect 42294 187954 42914 223398
rect 42294 187718 42326 187954
rect 42562 187718 42646 187954
rect 42882 187718 42914 187954
rect 42294 187634 42914 187718
rect 42294 187398 42326 187634
rect 42562 187398 42646 187634
rect 42882 187398 42914 187634
rect 42294 151954 42914 187398
rect 42294 151718 42326 151954
rect 42562 151718 42646 151954
rect 42882 151718 42914 151954
rect 42294 151634 42914 151718
rect 42294 151398 42326 151634
rect 42562 151398 42646 151634
rect 42882 151398 42914 151634
rect 42294 115954 42914 151398
rect 42294 115718 42326 115954
rect 42562 115718 42646 115954
rect 42882 115718 42914 115954
rect 42294 115634 42914 115718
rect 42294 115398 42326 115634
rect 42562 115398 42646 115634
rect 42882 115398 42914 115634
rect 42294 79954 42914 115398
rect 42294 79718 42326 79954
rect 42562 79718 42646 79954
rect 42882 79718 42914 79954
rect 42294 79634 42914 79718
rect 42294 79398 42326 79634
rect 42562 79398 42646 79634
rect 42882 79398 42914 79634
rect 42294 43954 42914 79398
rect 42294 43718 42326 43954
rect 42562 43718 42646 43954
rect 42882 43718 42914 43954
rect 42294 43634 42914 43718
rect 42294 43398 42326 43634
rect 42562 43398 42646 43634
rect 42882 43398 42914 43634
rect 42294 7954 42914 43398
rect 42294 7718 42326 7954
rect 42562 7718 42646 7954
rect 42882 7718 42914 7954
rect 42294 7634 42914 7718
rect 42294 7398 42326 7634
rect 42562 7398 42646 7634
rect 42882 7398 42914 7634
rect 42294 -1306 42914 7398
rect 42294 -1542 42326 -1306
rect 42562 -1542 42646 -1306
rect 42882 -1542 42914 -1306
rect 42294 -1626 42914 -1542
rect 42294 -1862 42326 -1626
rect 42562 -1862 42646 -1626
rect 42882 -1862 42914 -1626
rect 42294 -7654 42914 -1862
rect 46794 706758 47414 711590
rect 46794 706522 46826 706758
rect 47062 706522 47146 706758
rect 47382 706522 47414 706758
rect 46794 706438 47414 706522
rect 46794 706202 46826 706438
rect 47062 706202 47146 706438
rect 47382 706202 47414 706438
rect 46794 696454 47414 706202
rect 46794 696218 46826 696454
rect 47062 696218 47146 696454
rect 47382 696218 47414 696454
rect 46794 696134 47414 696218
rect 46794 695898 46826 696134
rect 47062 695898 47146 696134
rect 47382 695898 47414 696134
rect 46794 660454 47414 695898
rect 46794 660218 46826 660454
rect 47062 660218 47146 660454
rect 47382 660218 47414 660454
rect 46794 660134 47414 660218
rect 46794 659898 46826 660134
rect 47062 659898 47146 660134
rect 47382 659898 47414 660134
rect 46794 624454 47414 659898
rect 46794 624218 46826 624454
rect 47062 624218 47146 624454
rect 47382 624218 47414 624454
rect 46794 624134 47414 624218
rect 46794 623898 46826 624134
rect 47062 623898 47146 624134
rect 47382 623898 47414 624134
rect 46794 588454 47414 623898
rect 46794 588218 46826 588454
rect 47062 588218 47146 588454
rect 47382 588218 47414 588454
rect 46794 588134 47414 588218
rect 46794 587898 46826 588134
rect 47062 587898 47146 588134
rect 47382 587898 47414 588134
rect 46794 552454 47414 587898
rect 46794 552218 46826 552454
rect 47062 552218 47146 552454
rect 47382 552218 47414 552454
rect 46794 552134 47414 552218
rect 46794 551898 46826 552134
rect 47062 551898 47146 552134
rect 47382 551898 47414 552134
rect 46794 516454 47414 551898
rect 46794 516218 46826 516454
rect 47062 516218 47146 516454
rect 47382 516218 47414 516454
rect 46794 516134 47414 516218
rect 46794 515898 46826 516134
rect 47062 515898 47146 516134
rect 47382 515898 47414 516134
rect 46794 480454 47414 515898
rect 46794 480218 46826 480454
rect 47062 480218 47146 480454
rect 47382 480218 47414 480454
rect 46794 480134 47414 480218
rect 46794 479898 46826 480134
rect 47062 479898 47146 480134
rect 47382 479898 47414 480134
rect 46794 444454 47414 479898
rect 46794 444218 46826 444454
rect 47062 444218 47146 444454
rect 47382 444218 47414 444454
rect 46794 444134 47414 444218
rect 46794 443898 46826 444134
rect 47062 443898 47146 444134
rect 47382 443898 47414 444134
rect 46794 408454 47414 443898
rect 46794 408218 46826 408454
rect 47062 408218 47146 408454
rect 47382 408218 47414 408454
rect 46794 408134 47414 408218
rect 46794 407898 46826 408134
rect 47062 407898 47146 408134
rect 47382 407898 47414 408134
rect 46794 372454 47414 407898
rect 46794 372218 46826 372454
rect 47062 372218 47146 372454
rect 47382 372218 47414 372454
rect 46794 372134 47414 372218
rect 46794 371898 46826 372134
rect 47062 371898 47146 372134
rect 47382 371898 47414 372134
rect 46794 336454 47414 371898
rect 46794 336218 46826 336454
rect 47062 336218 47146 336454
rect 47382 336218 47414 336454
rect 46794 336134 47414 336218
rect 46794 335898 46826 336134
rect 47062 335898 47146 336134
rect 47382 335898 47414 336134
rect 46794 300454 47414 335898
rect 46794 300218 46826 300454
rect 47062 300218 47146 300454
rect 47382 300218 47414 300454
rect 46794 300134 47414 300218
rect 46794 299898 46826 300134
rect 47062 299898 47146 300134
rect 47382 299898 47414 300134
rect 46794 264454 47414 299898
rect 46794 264218 46826 264454
rect 47062 264218 47146 264454
rect 47382 264218 47414 264454
rect 46794 264134 47414 264218
rect 46794 263898 46826 264134
rect 47062 263898 47146 264134
rect 47382 263898 47414 264134
rect 46794 228454 47414 263898
rect 46794 228218 46826 228454
rect 47062 228218 47146 228454
rect 47382 228218 47414 228454
rect 46794 228134 47414 228218
rect 46794 227898 46826 228134
rect 47062 227898 47146 228134
rect 47382 227898 47414 228134
rect 46794 192454 47414 227898
rect 46794 192218 46826 192454
rect 47062 192218 47146 192454
rect 47382 192218 47414 192454
rect 46794 192134 47414 192218
rect 46794 191898 46826 192134
rect 47062 191898 47146 192134
rect 47382 191898 47414 192134
rect 46794 156454 47414 191898
rect 46794 156218 46826 156454
rect 47062 156218 47146 156454
rect 47382 156218 47414 156454
rect 46794 156134 47414 156218
rect 46794 155898 46826 156134
rect 47062 155898 47146 156134
rect 47382 155898 47414 156134
rect 46794 120454 47414 155898
rect 46794 120218 46826 120454
rect 47062 120218 47146 120454
rect 47382 120218 47414 120454
rect 46794 120134 47414 120218
rect 46794 119898 46826 120134
rect 47062 119898 47146 120134
rect 47382 119898 47414 120134
rect 46794 84454 47414 119898
rect 46794 84218 46826 84454
rect 47062 84218 47146 84454
rect 47382 84218 47414 84454
rect 46794 84134 47414 84218
rect 46794 83898 46826 84134
rect 47062 83898 47146 84134
rect 47382 83898 47414 84134
rect 46794 48454 47414 83898
rect 46794 48218 46826 48454
rect 47062 48218 47146 48454
rect 47382 48218 47414 48454
rect 46794 48134 47414 48218
rect 46794 47898 46826 48134
rect 47062 47898 47146 48134
rect 47382 47898 47414 48134
rect 46794 12454 47414 47898
rect 46794 12218 46826 12454
rect 47062 12218 47146 12454
rect 47382 12218 47414 12454
rect 46794 12134 47414 12218
rect 46794 11898 46826 12134
rect 47062 11898 47146 12134
rect 47382 11898 47414 12134
rect 46794 -2266 47414 11898
rect 46794 -2502 46826 -2266
rect 47062 -2502 47146 -2266
rect 47382 -2502 47414 -2266
rect 46794 -2586 47414 -2502
rect 46794 -2822 46826 -2586
rect 47062 -2822 47146 -2586
rect 47382 -2822 47414 -2586
rect 46794 -7654 47414 -2822
rect 51294 707718 51914 711590
rect 51294 707482 51326 707718
rect 51562 707482 51646 707718
rect 51882 707482 51914 707718
rect 51294 707398 51914 707482
rect 51294 707162 51326 707398
rect 51562 707162 51646 707398
rect 51882 707162 51914 707398
rect 51294 700954 51914 707162
rect 51294 700718 51326 700954
rect 51562 700718 51646 700954
rect 51882 700718 51914 700954
rect 51294 700634 51914 700718
rect 51294 700398 51326 700634
rect 51562 700398 51646 700634
rect 51882 700398 51914 700634
rect 51294 664954 51914 700398
rect 51294 664718 51326 664954
rect 51562 664718 51646 664954
rect 51882 664718 51914 664954
rect 51294 664634 51914 664718
rect 51294 664398 51326 664634
rect 51562 664398 51646 664634
rect 51882 664398 51914 664634
rect 51294 628954 51914 664398
rect 51294 628718 51326 628954
rect 51562 628718 51646 628954
rect 51882 628718 51914 628954
rect 51294 628634 51914 628718
rect 51294 628398 51326 628634
rect 51562 628398 51646 628634
rect 51882 628398 51914 628634
rect 51294 592954 51914 628398
rect 51294 592718 51326 592954
rect 51562 592718 51646 592954
rect 51882 592718 51914 592954
rect 51294 592634 51914 592718
rect 51294 592398 51326 592634
rect 51562 592398 51646 592634
rect 51882 592398 51914 592634
rect 51294 556954 51914 592398
rect 51294 556718 51326 556954
rect 51562 556718 51646 556954
rect 51882 556718 51914 556954
rect 51294 556634 51914 556718
rect 51294 556398 51326 556634
rect 51562 556398 51646 556634
rect 51882 556398 51914 556634
rect 51294 520954 51914 556398
rect 51294 520718 51326 520954
rect 51562 520718 51646 520954
rect 51882 520718 51914 520954
rect 51294 520634 51914 520718
rect 51294 520398 51326 520634
rect 51562 520398 51646 520634
rect 51882 520398 51914 520634
rect 51294 484954 51914 520398
rect 51294 484718 51326 484954
rect 51562 484718 51646 484954
rect 51882 484718 51914 484954
rect 51294 484634 51914 484718
rect 51294 484398 51326 484634
rect 51562 484398 51646 484634
rect 51882 484398 51914 484634
rect 51294 448954 51914 484398
rect 51294 448718 51326 448954
rect 51562 448718 51646 448954
rect 51882 448718 51914 448954
rect 51294 448634 51914 448718
rect 51294 448398 51326 448634
rect 51562 448398 51646 448634
rect 51882 448398 51914 448634
rect 51294 412954 51914 448398
rect 51294 412718 51326 412954
rect 51562 412718 51646 412954
rect 51882 412718 51914 412954
rect 51294 412634 51914 412718
rect 51294 412398 51326 412634
rect 51562 412398 51646 412634
rect 51882 412398 51914 412634
rect 51294 376954 51914 412398
rect 51294 376718 51326 376954
rect 51562 376718 51646 376954
rect 51882 376718 51914 376954
rect 51294 376634 51914 376718
rect 51294 376398 51326 376634
rect 51562 376398 51646 376634
rect 51882 376398 51914 376634
rect 51294 340954 51914 376398
rect 51294 340718 51326 340954
rect 51562 340718 51646 340954
rect 51882 340718 51914 340954
rect 51294 340634 51914 340718
rect 51294 340398 51326 340634
rect 51562 340398 51646 340634
rect 51882 340398 51914 340634
rect 51294 304954 51914 340398
rect 51294 304718 51326 304954
rect 51562 304718 51646 304954
rect 51882 304718 51914 304954
rect 51294 304634 51914 304718
rect 51294 304398 51326 304634
rect 51562 304398 51646 304634
rect 51882 304398 51914 304634
rect 51294 268954 51914 304398
rect 51294 268718 51326 268954
rect 51562 268718 51646 268954
rect 51882 268718 51914 268954
rect 51294 268634 51914 268718
rect 51294 268398 51326 268634
rect 51562 268398 51646 268634
rect 51882 268398 51914 268634
rect 51294 232954 51914 268398
rect 51294 232718 51326 232954
rect 51562 232718 51646 232954
rect 51882 232718 51914 232954
rect 51294 232634 51914 232718
rect 51294 232398 51326 232634
rect 51562 232398 51646 232634
rect 51882 232398 51914 232634
rect 51294 196954 51914 232398
rect 51294 196718 51326 196954
rect 51562 196718 51646 196954
rect 51882 196718 51914 196954
rect 51294 196634 51914 196718
rect 51294 196398 51326 196634
rect 51562 196398 51646 196634
rect 51882 196398 51914 196634
rect 51294 160954 51914 196398
rect 51294 160718 51326 160954
rect 51562 160718 51646 160954
rect 51882 160718 51914 160954
rect 51294 160634 51914 160718
rect 51294 160398 51326 160634
rect 51562 160398 51646 160634
rect 51882 160398 51914 160634
rect 51294 124954 51914 160398
rect 51294 124718 51326 124954
rect 51562 124718 51646 124954
rect 51882 124718 51914 124954
rect 51294 124634 51914 124718
rect 51294 124398 51326 124634
rect 51562 124398 51646 124634
rect 51882 124398 51914 124634
rect 51294 88954 51914 124398
rect 51294 88718 51326 88954
rect 51562 88718 51646 88954
rect 51882 88718 51914 88954
rect 51294 88634 51914 88718
rect 51294 88398 51326 88634
rect 51562 88398 51646 88634
rect 51882 88398 51914 88634
rect 51294 52954 51914 88398
rect 51294 52718 51326 52954
rect 51562 52718 51646 52954
rect 51882 52718 51914 52954
rect 51294 52634 51914 52718
rect 51294 52398 51326 52634
rect 51562 52398 51646 52634
rect 51882 52398 51914 52634
rect 51294 16954 51914 52398
rect 51294 16718 51326 16954
rect 51562 16718 51646 16954
rect 51882 16718 51914 16954
rect 51294 16634 51914 16718
rect 51294 16398 51326 16634
rect 51562 16398 51646 16634
rect 51882 16398 51914 16634
rect 51294 -3226 51914 16398
rect 51294 -3462 51326 -3226
rect 51562 -3462 51646 -3226
rect 51882 -3462 51914 -3226
rect 51294 -3546 51914 -3462
rect 51294 -3782 51326 -3546
rect 51562 -3782 51646 -3546
rect 51882 -3782 51914 -3546
rect 51294 -7654 51914 -3782
rect 55794 708678 56414 711590
rect 55794 708442 55826 708678
rect 56062 708442 56146 708678
rect 56382 708442 56414 708678
rect 55794 708358 56414 708442
rect 55794 708122 55826 708358
rect 56062 708122 56146 708358
rect 56382 708122 56414 708358
rect 55794 669454 56414 708122
rect 55794 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 56414 669454
rect 55794 669134 56414 669218
rect 55794 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 56414 669134
rect 55794 633454 56414 668898
rect 55794 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 56414 633454
rect 55794 633134 56414 633218
rect 55794 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 56414 633134
rect 55794 597454 56414 632898
rect 55794 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 56414 597454
rect 55794 597134 56414 597218
rect 55794 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 56414 597134
rect 55794 561454 56414 596898
rect 55794 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 56414 561454
rect 55794 561134 56414 561218
rect 55794 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 56414 561134
rect 55794 525454 56414 560898
rect 55794 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 56414 525454
rect 55794 525134 56414 525218
rect 55794 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 56414 525134
rect 55794 489454 56414 524898
rect 55794 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 56414 489454
rect 55794 489134 56414 489218
rect 55794 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 56414 489134
rect 55794 453454 56414 488898
rect 55794 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 56414 453454
rect 55794 453134 56414 453218
rect 55794 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 56414 453134
rect 55794 417454 56414 452898
rect 55794 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 56414 417454
rect 55794 417134 56414 417218
rect 55794 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 56414 417134
rect 55794 381454 56414 416898
rect 55794 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 56414 381454
rect 55794 381134 56414 381218
rect 55794 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 56414 381134
rect 55794 345454 56414 380898
rect 55794 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 56414 345454
rect 55794 345134 56414 345218
rect 55794 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 56414 345134
rect 55794 309454 56414 344898
rect 55794 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 56414 309454
rect 55794 309134 56414 309218
rect 55794 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 56414 309134
rect 55794 273454 56414 308898
rect 55794 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 56414 273454
rect 55794 273134 56414 273218
rect 55794 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 56414 273134
rect 55794 237454 56414 272898
rect 55794 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 56414 237454
rect 55794 237134 56414 237218
rect 55794 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 56414 237134
rect 55794 201454 56414 236898
rect 55794 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 56414 201454
rect 55794 201134 56414 201218
rect 55794 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 56414 201134
rect 55794 165454 56414 200898
rect 55794 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 56414 165454
rect 55794 165134 56414 165218
rect 55794 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 56414 165134
rect 55794 129454 56414 164898
rect 55794 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 56414 129454
rect 55794 129134 56414 129218
rect 55794 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 56414 129134
rect 55794 93454 56414 128898
rect 55794 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 56414 93454
rect 55794 93134 56414 93218
rect 55794 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 56414 93134
rect 55794 57454 56414 92898
rect 55794 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 56414 57454
rect 55794 57134 56414 57218
rect 55794 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 56414 57134
rect 55794 21454 56414 56898
rect 55794 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 56414 21454
rect 55794 21134 56414 21218
rect 55794 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 56414 21134
rect 55794 -4186 56414 20898
rect 55794 -4422 55826 -4186
rect 56062 -4422 56146 -4186
rect 56382 -4422 56414 -4186
rect 55794 -4506 56414 -4422
rect 55794 -4742 55826 -4506
rect 56062 -4742 56146 -4506
rect 56382 -4742 56414 -4506
rect 55794 -7654 56414 -4742
rect 60294 709638 60914 711590
rect 60294 709402 60326 709638
rect 60562 709402 60646 709638
rect 60882 709402 60914 709638
rect 60294 709318 60914 709402
rect 60294 709082 60326 709318
rect 60562 709082 60646 709318
rect 60882 709082 60914 709318
rect 60294 673954 60914 709082
rect 60294 673718 60326 673954
rect 60562 673718 60646 673954
rect 60882 673718 60914 673954
rect 60294 673634 60914 673718
rect 60294 673398 60326 673634
rect 60562 673398 60646 673634
rect 60882 673398 60914 673634
rect 60294 637954 60914 673398
rect 60294 637718 60326 637954
rect 60562 637718 60646 637954
rect 60882 637718 60914 637954
rect 60294 637634 60914 637718
rect 60294 637398 60326 637634
rect 60562 637398 60646 637634
rect 60882 637398 60914 637634
rect 60294 601954 60914 637398
rect 60294 601718 60326 601954
rect 60562 601718 60646 601954
rect 60882 601718 60914 601954
rect 60294 601634 60914 601718
rect 60294 601398 60326 601634
rect 60562 601398 60646 601634
rect 60882 601398 60914 601634
rect 60294 565954 60914 601398
rect 60294 565718 60326 565954
rect 60562 565718 60646 565954
rect 60882 565718 60914 565954
rect 60294 565634 60914 565718
rect 60294 565398 60326 565634
rect 60562 565398 60646 565634
rect 60882 565398 60914 565634
rect 60294 529954 60914 565398
rect 60294 529718 60326 529954
rect 60562 529718 60646 529954
rect 60882 529718 60914 529954
rect 60294 529634 60914 529718
rect 60294 529398 60326 529634
rect 60562 529398 60646 529634
rect 60882 529398 60914 529634
rect 60294 493954 60914 529398
rect 60294 493718 60326 493954
rect 60562 493718 60646 493954
rect 60882 493718 60914 493954
rect 60294 493634 60914 493718
rect 60294 493398 60326 493634
rect 60562 493398 60646 493634
rect 60882 493398 60914 493634
rect 60294 457954 60914 493398
rect 60294 457718 60326 457954
rect 60562 457718 60646 457954
rect 60882 457718 60914 457954
rect 60294 457634 60914 457718
rect 60294 457398 60326 457634
rect 60562 457398 60646 457634
rect 60882 457398 60914 457634
rect 60294 421954 60914 457398
rect 60294 421718 60326 421954
rect 60562 421718 60646 421954
rect 60882 421718 60914 421954
rect 60294 421634 60914 421718
rect 60294 421398 60326 421634
rect 60562 421398 60646 421634
rect 60882 421398 60914 421634
rect 60294 385954 60914 421398
rect 60294 385718 60326 385954
rect 60562 385718 60646 385954
rect 60882 385718 60914 385954
rect 60294 385634 60914 385718
rect 60294 385398 60326 385634
rect 60562 385398 60646 385634
rect 60882 385398 60914 385634
rect 60294 349954 60914 385398
rect 60294 349718 60326 349954
rect 60562 349718 60646 349954
rect 60882 349718 60914 349954
rect 60294 349634 60914 349718
rect 60294 349398 60326 349634
rect 60562 349398 60646 349634
rect 60882 349398 60914 349634
rect 60294 313954 60914 349398
rect 60294 313718 60326 313954
rect 60562 313718 60646 313954
rect 60882 313718 60914 313954
rect 60294 313634 60914 313718
rect 60294 313398 60326 313634
rect 60562 313398 60646 313634
rect 60882 313398 60914 313634
rect 60294 277954 60914 313398
rect 60294 277718 60326 277954
rect 60562 277718 60646 277954
rect 60882 277718 60914 277954
rect 60294 277634 60914 277718
rect 60294 277398 60326 277634
rect 60562 277398 60646 277634
rect 60882 277398 60914 277634
rect 60294 241954 60914 277398
rect 60294 241718 60326 241954
rect 60562 241718 60646 241954
rect 60882 241718 60914 241954
rect 60294 241634 60914 241718
rect 60294 241398 60326 241634
rect 60562 241398 60646 241634
rect 60882 241398 60914 241634
rect 60294 205954 60914 241398
rect 60294 205718 60326 205954
rect 60562 205718 60646 205954
rect 60882 205718 60914 205954
rect 60294 205634 60914 205718
rect 60294 205398 60326 205634
rect 60562 205398 60646 205634
rect 60882 205398 60914 205634
rect 60294 169954 60914 205398
rect 60294 169718 60326 169954
rect 60562 169718 60646 169954
rect 60882 169718 60914 169954
rect 60294 169634 60914 169718
rect 60294 169398 60326 169634
rect 60562 169398 60646 169634
rect 60882 169398 60914 169634
rect 60294 133954 60914 169398
rect 60294 133718 60326 133954
rect 60562 133718 60646 133954
rect 60882 133718 60914 133954
rect 60294 133634 60914 133718
rect 60294 133398 60326 133634
rect 60562 133398 60646 133634
rect 60882 133398 60914 133634
rect 60294 97954 60914 133398
rect 60294 97718 60326 97954
rect 60562 97718 60646 97954
rect 60882 97718 60914 97954
rect 60294 97634 60914 97718
rect 60294 97398 60326 97634
rect 60562 97398 60646 97634
rect 60882 97398 60914 97634
rect 60294 61954 60914 97398
rect 60294 61718 60326 61954
rect 60562 61718 60646 61954
rect 60882 61718 60914 61954
rect 60294 61634 60914 61718
rect 60294 61398 60326 61634
rect 60562 61398 60646 61634
rect 60882 61398 60914 61634
rect 60294 25954 60914 61398
rect 60294 25718 60326 25954
rect 60562 25718 60646 25954
rect 60882 25718 60914 25954
rect 60294 25634 60914 25718
rect 60294 25398 60326 25634
rect 60562 25398 60646 25634
rect 60882 25398 60914 25634
rect 60294 -5146 60914 25398
rect 60294 -5382 60326 -5146
rect 60562 -5382 60646 -5146
rect 60882 -5382 60914 -5146
rect 60294 -5466 60914 -5382
rect 60294 -5702 60326 -5466
rect 60562 -5702 60646 -5466
rect 60882 -5702 60914 -5466
rect 60294 -7654 60914 -5702
rect 64794 710598 65414 711590
rect 64794 710362 64826 710598
rect 65062 710362 65146 710598
rect 65382 710362 65414 710598
rect 64794 710278 65414 710362
rect 64794 710042 64826 710278
rect 65062 710042 65146 710278
rect 65382 710042 65414 710278
rect 64794 678454 65414 710042
rect 64794 678218 64826 678454
rect 65062 678218 65146 678454
rect 65382 678218 65414 678454
rect 64794 678134 65414 678218
rect 64794 677898 64826 678134
rect 65062 677898 65146 678134
rect 65382 677898 65414 678134
rect 64794 642454 65414 677898
rect 64794 642218 64826 642454
rect 65062 642218 65146 642454
rect 65382 642218 65414 642454
rect 64794 642134 65414 642218
rect 64794 641898 64826 642134
rect 65062 641898 65146 642134
rect 65382 641898 65414 642134
rect 64794 606454 65414 641898
rect 64794 606218 64826 606454
rect 65062 606218 65146 606454
rect 65382 606218 65414 606454
rect 64794 606134 65414 606218
rect 64794 605898 64826 606134
rect 65062 605898 65146 606134
rect 65382 605898 65414 606134
rect 64794 570454 65414 605898
rect 64794 570218 64826 570454
rect 65062 570218 65146 570454
rect 65382 570218 65414 570454
rect 64794 570134 65414 570218
rect 64794 569898 64826 570134
rect 65062 569898 65146 570134
rect 65382 569898 65414 570134
rect 64794 534454 65414 569898
rect 64794 534218 64826 534454
rect 65062 534218 65146 534454
rect 65382 534218 65414 534454
rect 64794 534134 65414 534218
rect 64794 533898 64826 534134
rect 65062 533898 65146 534134
rect 65382 533898 65414 534134
rect 64794 498454 65414 533898
rect 64794 498218 64826 498454
rect 65062 498218 65146 498454
rect 65382 498218 65414 498454
rect 64794 498134 65414 498218
rect 64794 497898 64826 498134
rect 65062 497898 65146 498134
rect 65382 497898 65414 498134
rect 64794 462454 65414 497898
rect 64794 462218 64826 462454
rect 65062 462218 65146 462454
rect 65382 462218 65414 462454
rect 64794 462134 65414 462218
rect 64794 461898 64826 462134
rect 65062 461898 65146 462134
rect 65382 461898 65414 462134
rect 64794 426454 65414 461898
rect 64794 426218 64826 426454
rect 65062 426218 65146 426454
rect 65382 426218 65414 426454
rect 64794 426134 65414 426218
rect 64794 425898 64826 426134
rect 65062 425898 65146 426134
rect 65382 425898 65414 426134
rect 64794 390454 65414 425898
rect 64794 390218 64826 390454
rect 65062 390218 65146 390454
rect 65382 390218 65414 390454
rect 64794 390134 65414 390218
rect 64794 389898 64826 390134
rect 65062 389898 65146 390134
rect 65382 389898 65414 390134
rect 64794 354454 65414 389898
rect 64794 354218 64826 354454
rect 65062 354218 65146 354454
rect 65382 354218 65414 354454
rect 64794 354134 65414 354218
rect 64794 353898 64826 354134
rect 65062 353898 65146 354134
rect 65382 353898 65414 354134
rect 64794 318454 65414 353898
rect 64794 318218 64826 318454
rect 65062 318218 65146 318454
rect 65382 318218 65414 318454
rect 64794 318134 65414 318218
rect 64794 317898 64826 318134
rect 65062 317898 65146 318134
rect 65382 317898 65414 318134
rect 64794 282454 65414 317898
rect 64794 282218 64826 282454
rect 65062 282218 65146 282454
rect 65382 282218 65414 282454
rect 64794 282134 65414 282218
rect 64794 281898 64826 282134
rect 65062 281898 65146 282134
rect 65382 281898 65414 282134
rect 64794 246454 65414 281898
rect 64794 246218 64826 246454
rect 65062 246218 65146 246454
rect 65382 246218 65414 246454
rect 64794 246134 65414 246218
rect 64794 245898 64826 246134
rect 65062 245898 65146 246134
rect 65382 245898 65414 246134
rect 64794 210454 65414 245898
rect 64794 210218 64826 210454
rect 65062 210218 65146 210454
rect 65382 210218 65414 210454
rect 64794 210134 65414 210218
rect 64794 209898 64826 210134
rect 65062 209898 65146 210134
rect 65382 209898 65414 210134
rect 64794 174454 65414 209898
rect 64794 174218 64826 174454
rect 65062 174218 65146 174454
rect 65382 174218 65414 174454
rect 64794 174134 65414 174218
rect 64794 173898 64826 174134
rect 65062 173898 65146 174134
rect 65382 173898 65414 174134
rect 64794 138454 65414 173898
rect 64794 138218 64826 138454
rect 65062 138218 65146 138454
rect 65382 138218 65414 138454
rect 64794 138134 65414 138218
rect 64794 137898 64826 138134
rect 65062 137898 65146 138134
rect 65382 137898 65414 138134
rect 64794 102454 65414 137898
rect 64794 102218 64826 102454
rect 65062 102218 65146 102454
rect 65382 102218 65414 102454
rect 64794 102134 65414 102218
rect 64794 101898 64826 102134
rect 65062 101898 65146 102134
rect 65382 101898 65414 102134
rect 64794 66454 65414 101898
rect 64794 66218 64826 66454
rect 65062 66218 65146 66454
rect 65382 66218 65414 66454
rect 64794 66134 65414 66218
rect 64794 65898 64826 66134
rect 65062 65898 65146 66134
rect 65382 65898 65414 66134
rect 64794 30454 65414 65898
rect 64794 30218 64826 30454
rect 65062 30218 65146 30454
rect 65382 30218 65414 30454
rect 64794 30134 65414 30218
rect 64794 29898 64826 30134
rect 65062 29898 65146 30134
rect 65382 29898 65414 30134
rect 64794 -6106 65414 29898
rect 64794 -6342 64826 -6106
rect 65062 -6342 65146 -6106
rect 65382 -6342 65414 -6106
rect 64794 -6426 65414 -6342
rect 64794 -6662 64826 -6426
rect 65062 -6662 65146 -6426
rect 65382 -6662 65414 -6426
rect 64794 -7654 65414 -6662
rect 69294 711558 69914 711590
rect 69294 711322 69326 711558
rect 69562 711322 69646 711558
rect 69882 711322 69914 711558
rect 69294 711238 69914 711322
rect 69294 711002 69326 711238
rect 69562 711002 69646 711238
rect 69882 711002 69914 711238
rect 69294 682954 69914 711002
rect 69294 682718 69326 682954
rect 69562 682718 69646 682954
rect 69882 682718 69914 682954
rect 69294 682634 69914 682718
rect 69294 682398 69326 682634
rect 69562 682398 69646 682634
rect 69882 682398 69914 682634
rect 69294 646954 69914 682398
rect 69294 646718 69326 646954
rect 69562 646718 69646 646954
rect 69882 646718 69914 646954
rect 69294 646634 69914 646718
rect 69294 646398 69326 646634
rect 69562 646398 69646 646634
rect 69882 646398 69914 646634
rect 69294 610954 69914 646398
rect 69294 610718 69326 610954
rect 69562 610718 69646 610954
rect 69882 610718 69914 610954
rect 69294 610634 69914 610718
rect 69294 610398 69326 610634
rect 69562 610398 69646 610634
rect 69882 610398 69914 610634
rect 69294 574954 69914 610398
rect 69294 574718 69326 574954
rect 69562 574718 69646 574954
rect 69882 574718 69914 574954
rect 69294 574634 69914 574718
rect 69294 574398 69326 574634
rect 69562 574398 69646 574634
rect 69882 574398 69914 574634
rect 69294 538954 69914 574398
rect 69294 538718 69326 538954
rect 69562 538718 69646 538954
rect 69882 538718 69914 538954
rect 69294 538634 69914 538718
rect 69294 538398 69326 538634
rect 69562 538398 69646 538634
rect 69882 538398 69914 538634
rect 69294 502954 69914 538398
rect 69294 502718 69326 502954
rect 69562 502718 69646 502954
rect 69882 502718 69914 502954
rect 69294 502634 69914 502718
rect 69294 502398 69326 502634
rect 69562 502398 69646 502634
rect 69882 502398 69914 502634
rect 69294 466954 69914 502398
rect 69294 466718 69326 466954
rect 69562 466718 69646 466954
rect 69882 466718 69914 466954
rect 69294 466634 69914 466718
rect 69294 466398 69326 466634
rect 69562 466398 69646 466634
rect 69882 466398 69914 466634
rect 69294 430954 69914 466398
rect 69294 430718 69326 430954
rect 69562 430718 69646 430954
rect 69882 430718 69914 430954
rect 69294 430634 69914 430718
rect 69294 430398 69326 430634
rect 69562 430398 69646 430634
rect 69882 430398 69914 430634
rect 69294 394954 69914 430398
rect 69294 394718 69326 394954
rect 69562 394718 69646 394954
rect 69882 394718 69914 394954
rect 69294 394634 69914 394718
rect 69294 394398 69326 394634
rect 69562 394398 69646 394634
rect 69882 394398 69914 394634
rect 69294 358954 69914 394398
rect 69294 358718 69326 358954
rect 69562 358718 69646 358954
rect 69882 358718 69914 358954
rect 69294 358634 69914 358718
rect 69294 358398 69326 358634
rect 69562 358398 69646 358634
rect 69882 358398 69914 358634
rect 69294 322954 69914 358398
rect 69294 322718 69326 322954
rect 69562 322718 69646 322954
rect 69882 322718 69914 322954
rect 69294 322634 69914 322718
rect 69294 322398 69326 322634
rect 69562 322398 69646 322634
rect 69882 322398 69914 322634
rect 69294 286954 69914 322398
rect 69294 286718 69326 286954
rect 69562 286718 69646 286954
rect 69882 286718 69914 286954
rect 69294 286634 69914 286718
rect 69294 286398 69326 286634
rect 69562 286398 69646 286634
rect 69882 286398 69914 286634
rect 69294 250954 69914 286398
rect 69294 250718 69326 250954
rect 69562 250718 69646 250954
rect 69882 250718 69914 250954
rect 69294 250634 69914 250718
rect 69294 250398 69326 250634
rect 69562 250398 69646 250634
rect 69882 250398 69914 250634
rect 69294 214954 69914 250398
rect 69294 214718 69326 214954
rect 69562 214718 69646 214954
rect 69882 214718 69914 214954
rect 69294 214634 69914 214718
rect 69294 214398 69326 214634
rect 69562 214398 69646 214634
rect 69882 214398 69914 214634
rect 69294 178954 69914 214398
rect 69294 178718 69326 178954
rect 69562 178718 69646 178954
rect 69882 178718 69914 178954
rect 69294 178634 69914 178718
rect 69294 178398 69326 178634
rect 69562 178398 69646 178634
rect 69882 178398 69914 178634
rect 69294 142954 69914 178398
rect 69294 142718 69326 142954
rect 69562 142718 69646 142954
rect 69882 142718 69914 142954
rect 69294 142634 69914 142718
rect 69294 142398 69326 142634
rect 69562 142398 69646 142634
rect 69882 142398 69914 142634
rect 69294 106954 69914 142398
rect 69294 106718 69326 106954
rect 69562 106718 69646 106954
rect 69882 106718 69914 106954
rect 69294 106634 69914 106718
rect 69294 106398 69326 106634
rect 69562 106398 69646 106634
rect 69882 106398 69914 106634
rect 69294 70954 69914 106398
rect 69294 70718 69326 70954
rect 69562 70718 69646 70954
rect 69882 70718 69914 70954
rect 69294 70634 69914 70718
rect 69294 70398 69326 70634
rect 69562 70398 69646 70634
rect 69882 70398 69914 70634
rect 69294 34954 69914 70398
rect 69294 34718 69326 34954
rect 69562 34718 69646 34954
rect 69882 34718 69914 34954
rect 69294 34634 69914 34718
rect 69294 34398 69326 34634
rect 69562 34398 69646 34634
rect 69882 34398 69914 34634
rect 69294 -7066 69914 34398
rect 69294 -7302 69326 -7066
rect 69562 -7302 69646 -7066
rect 69882 -7302 69914 -7066
rect 69294 -7386 69914 -7302
rect 69294 -7622 69326 -7386
rect 69562 -7622 69646 -7386
rect 69882 -7622 69914 -7386
rect 69294 -7654 69914 -7622
rect 73794 704838 74414 711590
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 73794 687454 74414 704282
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 651454 74414 686898
rect 73794 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 74414 651454
rect 73794 651134 74414 651218
rect 73794 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 74414 651134
rect 73794 615454 74414 650898
rect 73794 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 74414 615454
rect 73794 615134 74414 615218
rect 73794 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 74414 615134
rect 73794 579454 74414 614898
rect 73794 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 74414 579454
rect 73794 579134 74414 579218
rect 73794 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 74414 579134
rect 73794 543454 74414 578898
rect 73794 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 74414 543454
rect 73794 543134 74414 543218
rect 73794 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 74414 543134
rect 73794 507454 74414 542898
rect 73794 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 74414 507454
rect 73794 507134 74414 507218
rect 73794 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 74414 507134
rect 73794 471454 74414 506898
rect 73794 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 74414 471454
rect 73794 471134 74414 471218
rect 73794 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 74414 471134
rect 73794 435454 74414 470898
rect 73794 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 74414 435454
rect 73794 435134 74414 435218
rect 73794 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 74414 435134
rect 73794 399454 74414 434898
rect 73794 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 74414 399454
rect 73794 399134 74414 399218
rect 73794 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 74414 399134
rect 73794 363454 74414 398898
rect 73794 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 74414 363454
rect 73794 363134 74414 363218
rect 73794 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 74414 363134
rect 73794 327454 74414 362898
rect 73794 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 74414 327454
rect 73794 327134 74414 327218
rect 73794 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 74414 327134
rect 73794 291454 74414 326898
rect 73794 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 74414 291454
rect 73794 291134 74414 291218
rect 73794 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 74414 291134
rect 73794 255454 74414 290898
rect 73794 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 74414 255454
rect 73794 255134 74414 255218
rect 73794 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 74414 255134
rect 73794 219454 74414 254898
rect 73794 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 74414 219454
rect 73794 219134 74414 219218
rect 73794 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 74414 219134
rect 73794 183454 74414 218898
rect 73794 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 74414 183454
rect 73794 183134 74414 183218
rect 73794 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 74414 183134
rect 73794 147454 74414 182898
rect 73794 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 74414 147454
rect 73794 147134 74414 147218
rect 73794 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 74414 147134
rect 73794 111454 74414 146898
rect 73794 111218 73826 111454
rect 74062 111218 74146 111454
rect 74382 111218 74414 111454
rect 73794 111134 74414 111218
rect 73794 110898 73826 111134
rect 74062 110898 74146 111134
rect 74382 110898 74414 111134
rect 73794 75454 74414 110898
rect 73794 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 74414 75454
rect 73794 75134 74414 75218
rect 73794 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 74414 75134
rect 73794 39454 74414 74898
rect 73794 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 74414 39454
rect 73794 39134 74414 39218
rect 73794 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 74414 39134
rect 73794 3454 74414 38898
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -7654 74414 -902
rect 78294 705798 78914 711590
rect 78294 705562 78326 705798
rect 78562 705562 78646 705798
rect 78882 705562 78914 705798
rect 78294 705478 78914 705562
rect 78294 705242 78326 705478
rect 78562 705242 78646 705478
rect 78882 705242 78914 705478
rect 78294 691954 78914 705242
rect 78294 691718 78326 691954
rect 78562 691718 78646 691954
rect 78882 691718 78914 691954
rect 78294 691634 78914 691718
rect 78294 691398 78326 691634
rect 78562 691398 78646 691634
rect 78882 691398 78914 691634
rect 78294 655954 78914 691398
rect 78294 655718 78326 655954
rect 78562 655718 78646 655954
rect 78882 655718 78914 655954
rect 78294 655634 78914 655718
rect 78294 655398 78326 655634
rect 78562 655398 78646 655634
rect 78882 655398 78914 655634
rect 78294 619954 78914 655398
rect 78294 619718 78326 619954
rect 78562 619718 78646 619954
rect 78882 619718 78914 619954
rect 78294 619634 78914 619718
rect 78294 619398 78326 619634
rect 78562 619398 78646 619634
rect 78882 619398 78914 619634
rect 78294 583954 78914 619398
rect 78294 583718 78326 583954
rect 78562 583718 78646 583954
rect 78882 583718 78914 583954
rect 78294 583634 78914 583718
rect 78294 583398 78326 583634
rect 78562 583398 78646 583634
rect 78882 583398 78914 583634
rect 78294 547954 78914 583398
rect 78294 547718 78326 547954
rect 78562 547718 78646 547954
rect 78882 547718 78914 547954
rect 78294 547634 78914 547718
rect 78294 547398 78326 547634
rect 78562 547398 78646 547634
rect 78882 547398 78914 547634
rect 78294 511954 78914 547398
rect 78294 511718 78326 511954
rect 78562 511718 78646 511954
rect 78882 511718 78914 511954
rect 78294 511634 78914 511718
rect 78294 511398 78326 511634
rect 78562 511398 78646 511634
rect 78882 511398 78914 511634
rect 78294 475954 78914 511398
rect 78294 475718 78326 475954
rect 78562 475718 78646 475954
rect 78882 475718 78914 475954
rect 78294 475634 78914 475718
rect 78294 475398 78326 475634
rect 78562 475398 78646 475634
rect 78882 475398 78914 475634
rect 78294 439954 78914 475398
rect 78294 439718 78326 439954
rect 78562 439718 78646 439954
rect 78882 439718 78914 439954
rect 78294 439634 78914 439718
rect 78294 439398 78326 439634
rect 78562 439398 78646 439634
rect 78882 439398 78914 439634
rect 78294 403954 78914 439398
rect 78294 403718 78326 403954
rect 78562 403718 78646 403954
rect 78882 403718 78914 403954
rect 78294 403634 78914 403718
rect 78294 403398 78326 403634
rect 78562 403398 78646 403634
rect 78882 403398 78914 403634
rect 78294 367954 78914 403398
rect 78294 367718 78326 367954
rect 78562 367718 78646 367954
rect 78882 367718 78914 367954
rect 78294 367634 78914 367718
rect 78294 367398 78326 367634
rect 78562 367398 78646 367634
rect 78882 367398 78914 367634
rect 78294 331954 78914 367398
rect 78294 331718 78326 331954
rect 78562 331718 78646 331954
rect 78882 331718 78914 331954
rect 78294 331634 78914 331718
rect 78294 331398 78326 331634
rect 78562 331398 78646 331634
rect 78882 331398 78914 331634
rect 78294 295954 78914 331398
rect 78294 295718 78326 295954
rect 78562 295718 78646 295954
rect 78882 295718 78914 295954
rect 78294 295634 78914 295718
rect 78294 295398 78326 295634
rect 78562 295398 78646 295634
rect 78882 295398 78914 295634
rect 78294 259954 78914 295398
rect 78294 259718 78326 259954
rect 78562 259718 78646 259954
rect 78882 259718 78914 259954
rect 78294 259634 78914 259718
rect 78294 259398 78326 259634
rect 78562 259398 78646 259634
rect 78882 259398 78914 259634
rect 78294 223954 78914 259398
rect 78294 223718 78326 223954
rect 78562 223718 78646 223954
rect 78882 223718 78914 223954
rect 78294 223634 78914 223718
rect 78294 223398 78326 223634
rect 78562 223398 78646 223634
rect 78882 223398 78914 223634
rect 78294 187954 78914 223398
rect 78294 187718 78326 187954
rect 78562 187718 78646 187954
rect 78882 187718 78914 187954
rect 78294 187634 78914 187718
rect 78294 187398 78326 187634
rect 78562 187398 78646 187634
rect 78882 187398 78914 187634
rect 78294 151954 78914 187398
rect 78294 151718 78326 151954
rect 78562 151718 78646 151954
rect 78882 151718 78914 151954
rect 78294 151634 78914 151718
rect 78294 151398 78326 151634
rect 78562 151398 78646 151634
rect 78882 151398 78914 151634
rect 78294 115954 78914 151398
rect 78294 115718 78326 115954
rect 78562 115718 78646 115954
rect 78882 115718 78914 115954
rect 78294 115634 78914 115718
rect 78294 115398 78326 115634
rect 78562 115398 78646 115634
rect 78882 115398 78914 115634
rect 78294 79954 78914 115398
rect 78294 79718 78326 79954
rect 78562 79718 78646 79954
rect 78882 79718 78914 79954
rect 78294 79634 78914 79718
rect 78294 79398 78326 79634
rect 78562 79398 78646 79634
rect 78882 79398 78914 79634
rect 78294 43954 78914 79398
rect 78294 43718 78326 43954
rect 78562 43718 78646 43954
rect 78882 43718 78914 43954
rect 78294 43634 78914 43718
rect 78294 43398 78326 43634
rect 78562 43398 78646 43634
rect 78882 43398 78914 43634
rect 78294 7954 78914 43398
rect 78294 7718 78326 7954
rect 78562 7718 78646 7954
rect 78882 7718 78914 7954
rect 78294 7634 78914 7718
rect 78294 7398 78326 7634
rect 78562 7398 78646 7634
rect 78882 7398 78914 7634
rect 78294 -1306 78914 7398
rect 78294 -1542 78326 -1306
rect 78562 -1542 78646 -1306
rect 78882 -1542 78914 -1306
rect 78294 -1626 78914 -1542
rect 78294 -1862 78326 -1626
rect 78562 -1862 78646 -1626
rect 78882 -1862 78914 -1626
rect 78294 -7654 78914 -1862
rect 82794 706758 83414 711590
rect 82794 706522 82826 706758
rect 83062 706522 83146 706758
rect 83382 706522 83414 706758
rect 82794 706438 83414 706522
rect 82794 706202 82826 706438
rect 83062 706202 83146 706438
rect 83382 706202 83414 706438
rect 82794 696454 83414 706202
rect 82794 696218 82826 696454
rect 83062 696218 83146 696454
rect 83382 696218 83414 696454
rect 82794 696134 83414 696218
rect 82794 695898 82826 696134
rect 83062 695898 83146 696134
rect 83382 695898 83414 696134
rect 82794 660454 83414 695898
rect 82794 660218 82826 660454
rect 83062 660218 83146 660454
rect 83382 660218 83414 660454
rect 82794 660134 83414 660218
rect 82794 659898 82826 660134
rect 83062 659898 83146 660134
rect 83382 659898 83414 660134
rect 82794 624454 83414 659898
rect 82794 624218 82826 624454
rect 83062 624218 83146 624454
rect 83382 624218 83414 624454
rect 82794 624134 83414 624218
rect 82794 623898 82826 624134
rect 83062 623898 83146 624134
rect 83382 623898 83414 624134
rect 82794 588454 83414 623898
rect 82794 588218 82826 588454
rect 83062 588218 83146 588454
rect 83382 588218 83414 588454
rect 82794 588134 83414 588218
rect 82794 587898 82826 588134
rect 83062 587898 83146 588134
rect 83382 587898 83414 588134
rect 82794 552454 83414 587898
rect 82794 552218 82826 552454
rect 83062 552218 83146 552454
rect 83382 552218 83414 552454
rect 82794 552134 83414 552218
rect 82794 551898 82826 552134
rect 83062 551898 83146 552134
rect 83382 551898 83414 552134
rect 82794 516454 83414 551898
rect 82794 516218 82826 516454
rect 83062 516218 83146 516454
rect 83382 516218 83414 516454
rect 82794 516134 83414 516218
rect 82794 515898 82826 516134
rect 83062 515898 83146 516134
rect 83382 515898 83414 516134
rect 82794 480454 83414 515898
rect 82794 480218 82826 480454
rect 83062 480218 83146 480454
rect 83382 480218 83414 480454
rect 82794 480134 83414 480218
rect 82794 479898 82826 480134
rect 83062 479898 83146 480134
rect 83382 479898 83414 480134
rect 82794 444454 83414 479898
rect 82794 444218 82826 444454
rect 83062 444218 83146 444454
rect 83382 444218 83414 444454
rect 82794 444134 83414 444218
rect 82794 443898 82826 444134
rect 83062 443898 83146 444134
rect 83382 443898 83414 444134
rect 82794 408454 83414 443898
rect 82794 408218 82826 408454
rect 83062 408218 83146 408454
rect 83382 408218 83414 408454
rect 82794 408134 83414 408218
rect 82794 407898 82826 408134
rect 83062 407898 83146 408134
rect 83382 407898 83414 408134
rect 82794 372454 83414 407898
rect 82794 372218 82826 372454
rect 83062 372218 83146 372454
rect 83382 372218 83414 372454
rect 82794 372134 83414 372218
rect 82794 371898 82826 372134
rect 83062 371898 83146 372134
rect 83382 371898 83414 372134
rect 82794 336454 83414 371898
rect 82794 336218 82826 336454
rect 83062 336218 83146 336454
rect 83382 336218 83414 336454
rect 82794 336134 83414 336218
rect 82794 335898 82826 336134
rect 83062 335898 83146 336134
rect 83382 335898 83414 336134
rect 82794 300454 83414 335898
rect 82794 300218 82826 300454
rect 83062 300218 83146 300454
rect 83382 300218 83414 300454
rect 82794 300134 83414 300218
rect 82794 299898 82826 300134
rect 83062 299898 83146 300134
rect 83382 299898 83414 300134
rect 82794 264454 83414 299898
rect 82794 264218 82826 264454
rect 83062 264218 83146 264454
rect 83382 264218 83414 264454
rect 82794 264134 83414 264218
rect 82794 263898 82826 264134
rect 83062 263898 83146 264134
rect 83382 263898 83414 264134
rect 82794 228454 83414 263898
rect 82794 228218 82826 228454
rect 83062 228218 83146 228454
rect 83382 228218 83414 228454
rect 82794 228134 83414 228218
rect 82794 227898 82826 228134
rect 83062 227898 83146 228134
rect 83382 227898 83414 228134
rect 82794 192454 83414 227898
rect 82794 192218 82826 192454
rect 83062 192218 83146 192454
rect 83382 192218 83414 192454
rect 82794 192134 83414 192218
rect 82794 191898 82826 192134
rect 83062 191898 83146 192134
rect 83382 191898 83414 192134
rect 82794 156454 83414 191898
rect 82794 156218 82826 156454
rect 83062 156218 83146 156454
rect 83382 156218 83414 156454
rect 82794 156134 83414 156218
rect 82794 155898 82826 156134
rect 83062 155898 83146 156134
rect 83382 155898 83414 156134
rect 82794 120454 83414 155898
rect 82794 120218 82826 120454
rect 83062 120218 83146 120454
rect 83382 120218 83414 120454
rect 82794 120134 83414 120218
rect 82794 119898 82826 120134
rect 83062 119898 83146 120134
rect 83382 119898 83414 120134
rect 82794 84454 83414 119898
rect 82794 84218 82826 84454
rect 83062 84218 83146 84454
rect 83382 84218 83414 84454
rect 82794 84134 83414 84218
rect 82794 83898 82826 84134
rect 83062 83898 83146 84134
rect 83382 83898 83414 84134
rect 82794 48454 83414 83898
rect 82794 48218 82826 48454
rect 83062 48218 83146 48454
rect 83382 48218 83414 48454
rect 82794 48134 83414 48218
rect 82794 47898 82826 48134
rect 83062 47898 83146 48134
rect 83382 47898 83414 48134
rect 82794 12454 83414 47898
rect 82794 12218 82826 12454
rect 83062 12218 83146 12454
rect 83382 12218 83414 12454
rect 82794 12134 83414 12218
rect 82794 11898 82826 12134
rect 83062 11898 83146 12134
rect 83382 11898 83414 12134
rect 82794 -2266 83414 11898
rect 82794 -2502 82826 -2266
rect 83062 -2502 83146 -2266
rect 83382 -2502 83414 -2266
rect 82794 -2586 83414 -2502
rect 82794 -2822 82826 -2586
rect 83062 -2822 83146 -2586
rect 83382 -2822 83414 -2586
rect 82794 -7654 83414 -2822
rect 87294 707718 87914 711590
rect 87294 707482 87326 707718
rect 87562 707482 87646 707718
rect 87882 707482 87914 707718
rect 87294 707398 87914 707482
rect 87294 707162 87326 707398
rect 87562 707162 87646 707398
rect 87882 707162 87914 707398
rect 87294 700954 87914 707162
rect 87294 700718 87326 700954
rect 87562 700718 87646 700954
rect 87882 700718 87914 700954
rect 87294 700634 87914 700718
rect 87294 700398 87326 700634
rect 87562 700398 87646 700634
rect 87882 700398 87914 700634
rect 87294 664954 87914 700398
rect 87294 664718 87326 664954
rect 87562 664718 87646 664954
rect 87882 664718 87914 664954
rect 87294 664634 87914 664718
rect 87294 664398 87326 664634
rect 87562 664398 87646 664634
rect 87882 664398 87914 664634
rect 87294 628954 87914 664398
rect 87294 628718 87326 628954
rect 87562 628718 87646 628954
rect 87882 628718 87914 628954
rect 87294 628634 87914 628718
rect 87294 628398 87326 628634
rect 87562 628398 87646 628634
rect 87882 628398 87914 628634
rect 87294 592954 87914 628398
rect 87294 592718 87326 592954
rect 87562 592718 87646 592954
rect 87882 592718 87914 592954
rect 87294 592634 87914 592718
rect 87294 592398 87326 592634
rect 87562 592398 87646 592634
rect 87882 592398 87914 592634
rect 87294 556954 87914 592398
rect 87294 556718 87326 556954
rect 87562 556718 87646 556954
rect 87882 556718 87914 556954
rect 87294 556634 87914 556718
rect 87294 556398 87326 556634
rect 87562 556398 87646 556634
rect 87882 556398 87914 556634
rect 87294 520954 87914 556398
rect 87294 520718 87326 520954
rect 87562 520718 87646 520954
rect 87882 520718 87914 520954
rect 87294 520634 87914 520718
rect 87294 520398 87326 520634
rect 87562 520398 87646 520634
rect 87882 520398 87914 520634
rect 87294 484954 87914 520398
rect 87294 484718 87326 484954
rect 87562 484718 87646 484954
rect 87882 484718 87914 484954
rect 87294 484634 87914 484718
rect 87294 484398 87326 484634
rect 87562 484398 87646 484634
rect 87882 484398 87914 484634
rect 87294 448954 87914 484398
rect 87294 448718 87326 448954
rect 87562 448718 87646 448954
rect 87882 448718 87914 448954
rect 87294 448634 87914 448718
rect 87294 448398 87326 448634
rect 87562 448398 87646 448634
rect 87882 448398 87914 448634
rect 87294 412954 87914 448398
rect 87294 412718 87326 412954
rect 87562 412718 87646 412954
rect 87882 412718 87914 412954
rect 87294 412634 87914 412718
rect 87294 412398 87326 412634
rect 87562 412398 87646 412634
rect 87882 412398 87914 412634
rect 87294 376954 87914 412398
rect 87294 376718 87326 376954
rect 87562 376718 87646 376954
rect 87882 376718 87914 376954
rect 87294 376634 87914 376718
rect 87294 376398 87326 376634
rect 87562 376398 87646 376634
rect 87882 376398 87914 376634
rect 87294 340954 87914 376398
rect 87294 340718 87326 340954
rect 87562 340718 87646 340954
rect 87882 340718 87914 340954
rect 87294 340634 87914 340718
rect 87294 340398 87326 340634
rect 87562 340398 87646 340634
rect 87882 340398 87914 340634
rect 87294 304954 87914 340398
rect 87294 304718 87326 304954
rect 87562 304718 87646 304954
rect 87882 304718 87914 304954
rect 87294 304634 87914 304718
rect 87294 304398 87326 304634
rect 87562 304398 87646 304634
rect 87882 304398 87914 304634
rect 87294 268954 87914 304398
rect 87294 268718 87326 268954
rect 87562 268718 87646 268954
rect 87882 268718 87914 268954
rect 87294 268634 87914 268718
rect 87294 268398 87326 268634
rect 87562 268398 87646 268634
rect 87882 268398 87914 268634
rect 87294 232954 87914 268398
rect 87294 232718 87326 232954
rect 87562 232718 87646 232954
rect 87882 232718 87914 232954
rect 87294 232634 87914 232718
rect 87294 232398 87326 232634
rect 87562 232398 87646 232634
rect 87882 232398 87914 232634
rect 87294 196954 87914 232398
rect 87294 196718 87326 196954
rect 87562 196718 87646 196954
rect 87882 196718 87914 196954
rect 87294 196634 87914 196718
rect 87294 196398 87326 196634
rect 87562 196398 87646 196634
rect 87882 196398 87914 196634
rect 87294 160954 87914 196398
rect 87294 160718 87326 160954
rect 87562 160718 87646 160954
rect 87882 160718 87914 160954
rect 87294 160634 87914 160718
rect 87294 160398 87326 160634
rect 87562 160398 87646 160634
rect 87882 160398 87914 160634
rect 87294 124954 87914 160398
rect 87294 124718 87326 124954
rect 87562 124718 87646 124954
rect 87882 124718 87914 124954
rect 87294 124634 87914 124718
rect 87294 124398 87326 124634
rect 87562 124398 87646 124634
rect 87882 124398 87914 124634
rect 87294 88954 87914 124398
rect 87294 88718 87326 88954
rect 87562 88718 87646 88954
rect 87882 88718 87914 88954
rect 87294 88634 87914 88718
rect 87294 88398 87326 88634
rect 87562 88398 87646 88634
rect 87882 88398 87914 88634
rect 87294 52954 87914 88398
rect 87294 52718 87326 52954
rect 87562 52718 87646 52954
rect 87882 52718 87914 52954
rect 87294 52634 87914 52718
rect 87294 52398 87326 52634
rect 87562 52398 87646 52634
rect 87882 52398 87914 52634
rect 87294 16954 87914 52398
rect 87294 16718 87326 16954
rect 87562 16718 87646 16954
rect 87882 16718 87914 16954
rect 87294 16634 87914 16718
rect 87294 16398 87326 16634
rect 87562 16398 87646 16634
rect 87882 16398 87914 16634
rect 87294 -3226 87914 16398
rect 87294 -3462 87326 -3226
rect 87562 -3462 87646 -3226
rect 87882 -3462 87914 -3226
rect 87294 -3546 87914 -3462
rect 87294 -3782 87326 -3546
rect 87562 -3782 87646 -3546
rect 87882 -3782 87914 -3546
rect 87294 -7654 87914 -3782
rect 91794 708678 92414 711590
rect 91794 708442 91826 708678
rect 92062 708442 92146 708678
rect 92382 708442 92414 708678
rect 91794 708358 92414 708442
rect 91794 708122 91826 708358
rect 92062 708122 92146 708358
rect 92382 708122 92414 708358
rect 91794 669454 92414 708122
rect 91794 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 92414 669454
rect 91794 669134 92414 669218
rect 91794 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 92414 669134
rect 91794 633454 92414 668898
rect 91794 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 92414 633454
rect 91794 633134 92414 633218
rect 91794 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 92414 633134
rect 91794 597454 92414 632898
rect 91794 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 92414 597454
rect 91794 597134 92414 597218
rect 91794 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 92414 597134
rect 91794 561454 92414 596898
rect 91794 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 92414 561454
rect 91794 561134 92414 561218
rect 91794 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 92414 561134
rect 91794 525454 92414 560898
rect 91794 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 92414 525454
rect 91794 525134 92414 525218
rect 91794 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 92414 525134
rect 91794 489454 92414 524898
rect 91794 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 92414 489454
rect 91794 489134 92414 489218
rect 91794 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 92414 489134
rect 91794 453454 92414 488898
rect 91794 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 92414 453454
rect 91794 453134 92414 453218
rect 91794 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 92414 453134
rect 91794 417454 92414 452898
rect 91794 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 92414 417454
rect 91794 417134 92414 417218
rect 91794 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 92414 417134
rect 91794 381454 92414 416898
rect 91794 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 92414 381454
rect 91794 381134 92414 381218
rect 91794 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 92414 381134
rect 91794 345454 92414 380898
rect 91794 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 92414 345454
rect 91794 345134 92414 345218
rect 91794 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 92414 345134
rect 91794 309454 92414 344898
rect 91794 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 92414 309454
rect 91794 309134 92414 309218
rect 91794 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 92414 309134
rect 91794 273454 92414 308898
rect 91794 273218 91826 273454
rect 92062 273218 92146 273454
rect 92382 273218 92414 273454
rect 91794 273134 92414 273218
rect 91794 272898 91826 273134
rect 92062 272898 92146 273134
rect 92382 272898 92414 273134
rect 91794 237454 92414 272898
rect 91794 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 92414 237454
rect 91794 237134 92414 237218
rect 91794 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 92414 237134
rect 91794 201454 92414 236898
rect 91794 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 92414 201454
rect 91794 201134 92414 201218
rect 91794 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 92414 201134
rect 91794 165454 92414 200898
rect 91794 165218 91826 165454
rect 92062 165218 92146 165454
rect 92382 165218 92414 165454
rect 91794 165134 92414 165218
rect 91794 164898 91826 165134
rect 92062 164898 92146 165134
rect 92382 164898 92414 165134
rect 91794 129454 92414 164898
rect 91794 129218 91826 129454
rect 92062 129218 92146 129454
rect 92382 129218 92414 129454
rect 91794 129134 92414 129218
rect 91794 128898 91826 129134
rect 92062 128898 92146 129134
rect 92382 128898 92414 129134
rect 91794 93454 92414 128898
rect 91794 93218 91826 93454
rect 92062 93218 92146 93454
rect 92382 93218 92414 93454
rect 91794 93134 92414 93218
rect 91794 92898 91826 93134
rect 92062 92898 92146 93134
rect 92382 92898 92414 93134
rect 91794 57454 92414 92898
rect 91794 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 92414 57454
rect 91794 57134 92414 57218
rect 91794 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 92414 57134
rect 91794 21454 92414 56898
rect 91794 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 92414 21454
rect 91794 21134 92414 21218
rect 91794 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 92414 21134
rect 91794 -4186 92414 20898
rect 91794 -4422 91826 -4186
rect 92062 -4422 92146 -4186
rect 92382 -4422 92414 -4186
rect 91794 -4506 92414 -4422
rect 91794 -4742 91826 -4506
rect 92062 -4742 92146 -4506
rect 92382 -4742 92414 -4506
rect 91794 -7654 92414 -4742
rect 96294 709638 96914 711590
rect 96294 709402 96326 709638
rect 96562 709402 96646 709638
rect 96882 709402 96914 709638
rect 96294 709318 96914 709402
rect 96294 709082 96326 709318
rect 96562 709082 96646 709318
rect 96882 709082 96914 709318
rect 96294 673954 96914 709082
rect 96294 673718 96326 673954
rect 96562 673718 96646 673954
rect 96882 673718 96914 673954
rect 96294 673634 96914 673718
rect 96294 673398 96326 673634
rect 96562 673398 96646 673634
rect 96882 673398 96914 673634
rect 96294 637954 96914 673398
rect 96294 637718 96326 637954
rect 96562 637718 96646 637954
rect 96882 637718 96914 637954
rect 96294 637634 96914 637718
rect 96294 637398 96326 637634
rect 96562 637398 96646 637634
rect 96882 637398 96914 637634
rect 96294 601954 96914 637398
rect 96294 601718 96326 601954
rect 96562 601718 96646 601954
rect 96882 601718 96914 601954
rect 96294 601634 96914 601718
rect 96294 601398 96326 601634
rect 96562 601398 96646 601634
rect 96882 601398 96914 601634
rect 96294 565954 96914 601398
rect 100794 710598 101414 711590
rect 100794 710362 100826 710598
rect 101062 710362 101146 710598
rect 101382 710362 101414 710598
rect 100794 710278 101414 710362
rect 100794 710042 100826 710278
rect 101062 710042 101146 710278
rect 101382 710042 101414 710278
rect 100794 678454 101414 710042
rect 100794 678218 100826 678454
rect 101062 678218 101146 678454
rect 101382 678218 101414 678454
rect 100794 678134 101414 678218
rect 100794 677898 100826 678134
rect 101062 677898 101146 678134
rect 101382 677898 101414 678134
rect 100794 642454 101414 677898
rect 100794 642218 100826 642454
rect 101062 642218 101146 642454
rect 101382 642218 101414 642454
rect 100794 642134 101414 642218
rect 100794 641898 100826 642134
rect 101062 641898 101146 642134
rect 101382 641898 101414 642134
rect 100794 606454 101414 641898
rect 100794 606218 100826 606454
rect 101062 606218 101146 606454
rect 101382 606218 101414 606454
rect 100794 606134 101414 606218
rect 100794 605898 100826 606134
rect 101062 605898 101146 606134
rect 101382 605898 101414 606134
rect 100794 591292 101414 605898
rect 105294 711558 105914 711590
rect 105294 711322 105326 711558
rect 105562 711322 105646 711558
rect 105882 711322 105914 711558
rect 105294 711238 105914 711322
rect 105294 711002 105326 711238
rect 105562 711002 105646 711238
rect 105882 711002 105914 711238
rect 105294 682954 105914 711002
rect 105294 682718 105326 682954
rect 105562 682718 105646 682954
rect 105882 682718 105914 682954
rect 105294 682634 105914 682718
rect 105294 682398 105326 682634
rect 105562 682398 105646 682634
rect 105882 682398 105914 682634
rect 105294 646954 105914 682398
rect 105294 646718 105326 646954
rect 105562 646718 105646 646954
rect 105882 646718 105914 646954
rect 105294 646634 105914 646718
rect 105294 646398 105326 646634
rect 105562 646398 105646 646634
rect 105882 646398 105914 646634
rect 105294 610954 105914 646398
rect 105294 610718 105326 610954
rect 105562 610718 105646 610954
rect 105882 610718 105914 610954
rect 105294 610634 105914 610718
rect 105294 610398 105326 610634
rect 105562 610398 105646 610634
rect 105882 610398 105914 610634
rect 105294 591292 105914 610398
rect 109794 704838 110414 711590
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 687454 110414 704282
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 651454 110414 686898
rect 109794 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 110414 651454
rect 109794 651134 110414 651218
rect 109794 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 110414 651134
rect 109794 615454 110414 650898
rect 109794 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 110414 615454
rect 109794 615134 110414 615218
rect 109794 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 110414 615134
rect 109794 591292 110414 614898
rect 114294 705798 114914 711590
rect 114294 705562 114326 705798
rect 114562 705562 114646 705798
rect 114882 705562 114914 705798
rect 114294 705478 114914 705562
rect 114294 705242 114326 705478
rect 114562 705242 114646 705478
rect 114882 705242 114914 705478
rect 114294 691954 114914 705242
rect 114294 691718 114326 691954
rect 114562 691718 114646 691954
rect 114882 691718 114914 691954
rect 114294 691634 114914 691718
rect 114294 691398 114326 691634
rect 114562 691398 114646 691634
rect 114882 691398 114914 691634
rect 114294 655954 114914 691398
rect 114294 655718 114326 655954
rect 114562 655718 114646 655954
rect 114882 655718 114914 655954
rect 114294 655634 114914 655718
rect 114294 655398 114326 655634
rect 114562 655398 114646 655634
rect 114882 655398 114914 655634
rect 114294 619954 114914 655398
rect 114294 619718 114326 619954
rect 114562 619718 114646 619954
rect 114882 619718 114914 619954
rect 114294 619634 114914 619718
rect 114294 619398 114326 619634
rect 114562 619398 114646 619634
rect 114882 619398 114914 619634
rect 114294 591292 114914 619398
rect 118794 706758 119414 711590
rect 118794 706522 118826 706758
rect 119062 706522 119146 706758
rect 119382 706522 119414 706758
rect 118794 706438 119414 706522
rect 118794 706202 118826 706438
rect 119062 706202 119146 706438
rect 119382 706202 119414 706438
rect 118794 696454 119414 706202
rect 118794 696218 118826 696454
rect 119062 696218 119146 696454
rect 119382 696218 119414 696454
rect 118794 696134 119414 696218
rect 118794 695898 118826 696134
rect 119062 695898 119146 696134
rect 119382 695898 119414 696134
rect 118794 660454 119414 695898
rect 118794 660218 118826 660454
rect 119062 660218 119146 660454
rect 119382 660218 119414 660454
rect 118794 660134 119414 660218
rect 118794 659898 118826 660134
rect 119062 659898 119146 660134
rect 119382 659898 119414 660134
rect 118794 624454 119414 659898
rect 118794 624218 118826 624454
rect 119062 624218 119146 624454
rect 119382 624218 119414 624454
rect 118794 624134 119414 624218
rect 118794 623898 118826 624134
rect 119062 623898 119146 624134
rect 119382 623898 119414 624134
rect 118794 591292 119414 623898
rect 123294 707718 123914 711590
rect 123294 707482 123326 707718
rect 123562 707482 123646 707718
rect 123882 707482 123914 707718
rect 123294 707398 123914 707482
rect 123294 707162 123326 707398
rect 123562 707162 123646 707398
rect 123882 707162 123914 707398
rect 123294 700954 123914 707162
rect 123294 700718 123326 700954
rect 123562 700718 123646 700954
rect 123882 700718 123914 700954
rect 123294 700634 123914 700718
rect 123294 700398 123326 700634
rect 123562 700398 123646 700634
rect 123882 700398 123914 700634
rect 123294 664954 123914 700398
rect 123294 664718 123326 664954
rect 123562 664718 123646 664954
rect 123882 664718 123914 664954
rect 123294 664634 123914 664718
rect 123294 664398 123326 664634
rect 123562 664398 123646 664634
rect 123882 664398 123914 664634
rect 123294 628954 123914 664398
rect 123294 628718 123326 628954
rect 123562 628718 123646 628954
rect 123882 628718 123914 628954
rect 123294 628634 123914 628718
rect 123294 628398 123326 628634
rect 123562 628398 123646 628634
rect 123882 628398 123914 628634
rect 123294 592954 123914 628398
rect 123294 592718 123326 592954
rect 123562 592718 123646 592954
rect 123882 592718 123914 592954
rect 123294 592634 123914 592718
rect 123294 592398 123326 592634
rect 123562 592398 123646 592634
rect 123882 592398 123914 592634
rect 123294 591292 123914 592398
rect 127794 708678 128414 711590
rect 127794 708442 127826 708678
rect 128062 708442 128146 708678
rect 128382 708442 128414 708678
rect 127794 708358 128414 708442
rect 127794 708122 127826 708358
rect 128062 708122 128146 708358
rect 128382 708122 128414 708358
rect 127794 669454 128414 708122
rect 127794 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 128414 669454
rect 127794 669134 128414 669218
rect 127794 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 128414 669134
rect 127794 633454 128414 668898
rect 127794 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 128414 633454
rect 127794 633134 128414 633218
rect 127794 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 128414 633134
rect 127794 597454 128414 632898
rect 127794 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 128414 597454
rect 127794 597134 128414 597218
rect 127794 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 128414 597134
rect 127794 591292 128414 596898
rect 132294 709638 132914 711590
rect 132294 709402 132326 709638
rect 132562 709402 132646 709638
rect 132882 709402 132914 709638
rect 132294 709318 132914 709402
rect 132294 709082 132326 709318
rect 132562 709082 132646 709318
rect 132882 709082 132914 709318
rect 132294 673954 132914 709082
rect 132294 673718 132326 673954
rect 132562 673718 132646 673954
rect 132882 673718 132914 673954
rect 132294 673634 132914 673718
rect 132294 673398 132326 673634
rect 132562 673398 132646 673634
rect 132882 673398 132914 673634
rect 132294 637954 132914 673398
rect 132294 637718 132326 637954
rect 132562 637718 132646 637954
rect 132882 637718 132914 637954
rect 132294 637634 132914 637718
rect 132294 637398 132326 637634
rect 132562 637398 132646 637634
rect 132882 637398 132914 637634
rect 132294 601954 132914 637398
rect 132294 601718 132326 601954
rect 132562 601718 132646 601954
rect 132882 601718 132914 601954
rect 132294 601634 132914 601718
rect 132294 601398 132326 601634
rect 132562 601398 132646 601634
rect 132882 601398 132914 601634
rect 132294 591292 132914 601398
rect 136794 710598 137414 711590
rect 136794 710362 136826 710598
rect 137062 710362 137146 710598
rect 137382 710362 137414 710598
rect 136794 710278 137414 710362
rect 136794 710042 136826 710278
rect 137062 710042 137146 710278
rect 137382 710042 137414 710278
rect 136794 678454 137414 710042
rect 136794 678218 136826 678454
rect 137062 678218 137146 678454
rect 137382 678218 137414 678454
rect 136794 678134 137414 678218
rect 136794 677898 136826 678134
rect 137062 677898 137146 678134
rect 137382 677898 137414 678134
rect 136794 642454 137414 677898
rect 136794 642218 136826 642454
rect 137062 642218 137146 642454
rect 137382 642218 137414 642454
rect 136794 642134 137414 642218
rect 136794 641898 136826 642134
rect 137062 641898 137146 642134
rect 137382 641898 137414 642134
rect 136794 606454 137414 641898
rect 136794 606218 136826 606454
rect 137062 606218 137146 606454
rect 137382 606218 137414 606454
rect 136794 606134 137414 606218
rect 136794 605898 136826 606134
rect 137062 605898 137146 606134
rect 137382 605898 137414 606134
rect 136794 591292 137414 605898
rect 141294 711558 141914 711590
rect 141294 711322 141326 711558
rect 141562 711322 141646 711558
rect 141882 711322 141914 711558
rect 141294 711238 141914 711322
rect 141294 711002 141326 711238
rect 141562 711002 141646 711238
rect 141882 711002 141914 711238
rect 141294 682954 141914 711002
rect 141294 682718 141326 682954
rect 141562 682718 141646 682954
rect 141882 682718 141914 682954
rect 141294 682634 141914 682718
rect 141294 682398 141326 682634
rect 141562 682398 141646 682634
rect 141882 682398 141914 682634
rect 141294 646954 141914 682398
rect 141294 646718 141326 646954
rect 141562 646718 141646 646954
rect 141882 646718 141914 646954
rect 141294 646634 141914 646718
rect 141294 646398 141326 646634
rect 141562 646398 141646 646634
rect 141882 646398 141914 646634
rect 141294 610954 141914 646398
rect 141294 610718 141326 610954
rect 141562 610718 141646 610954
rect 141882 610718 141914 610954
rect 141294 610634 141914 610718
rect 141294 610398 141326 610634
rect 141562 610398 141646 610634
rect 141882 610398 141914 610634
rect 141294 591292 141914 610398
rect 145794 704838 146414 711590
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 687454 146414 704282
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 651454 146414 686898
rect 145794 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 146414 651454
rect 145794 651134 146414 651218
rect 145794 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 146414 651134
rect 145794 615454 146414 650898
rect 145794 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 146414 615454
rect 145794 615134 146414 615218
rect 145794 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 146414 615134
rect 145794 591292 146414 614898
rect 150294 705798 150914 711590
rect 150294 705562 150326 705798
rect 150562 705562 150646 705798
rect 150882 705562 150914 705798
rect 150294 705478 150914 705562
rect 150294 705242 150326 705478
rect 150562 705242 150646 705478
rect 150882 705242 150914 705478
rect 150294 691954 150914 705242
rect 150294 691718 150326 691954
rect 150562 691718 150646 691954
rect 150882 691718 150914 691954
rect 150294 691634 150914 691718
rect 150294 691398 150326 691634
rect 150562 691398 150646 691634
rect 150882 691398 150914 691634
rect 150294 655954 150914 691398
rect 150294 655718 150326 655954
rect 150562 655718 150646 655954
rect 150882 655718 150914 655954
rect 150294 655634 150914 655718
rect 150294 655398 150326 655634
rect 150562 655398 150646 655634
rect 150882 655398 150914 655634
rect 150294 619954 150914 655398
rect 150294 619718 150326 619954
rect 150562 619718 150646 619954
rect 150882 619718 150914 619954
rect 150294 619634 150914 619718
rect 150294 619398 150326 619634
rect 150562 619398 150646 619634
rect 150882 619398 150914 619634
rect 150294 591292 150914 619398
rect 154794 706758 155414 711590
rect 154794 706522 154826 706758
rect 155062 706522 155146 706758
rect 155382 706522 155414 706758
rect 154794 706438 155414 706522
rect 154794 706202 154826 706438
rect 155062 706202 155146 706438
rect 155382 706202 155414 706438
rect 154794 696454 155414 706202
rect 154794 696218 154826 696454
rect 155062 696218 155146 696454
rect 155382 696218 155414 696454
rect 154794 696134 155414 696218
rect 154794 695898 154826 696134
rect 155062 695898 155146 696134
rect 155382 695898 155414 696134
rect 154794 660454 155414 695898
rect 154794 660218 154826 660454
rect 155062 660218 155146 660454
rect 155382 660218 155414 660454
rect 154794 660134 155414 660218
rect 154794 659898 154826 660134
rect 155062 659898 155146 660134
rect 155382 659898 155414 660134
rect 154794 624454 155414 659898
rect 154794 624218 154826 624454
rect 155062 624218 155146 624454
rect 155382 624218 155414 624454
rect 154794 624134 155414 624218
rect 154794 623898 154826 624134
rect 155062 623898 155146 624134
rect 155382 623898 155414 624134
rect 154794 591292 155414 623898
rect 159294 707718 159914 711590
rect 159294 707482 159326 707718
rect 159562 707482 159646 707718
rect 159882 707482 159914 707718
rect 159294 707398 159914 707482
rect 159294 707162 159326 707398
rect 159562 707162 159646 707398
rect 159882 707162 159914 707398
rect 159294 700954 159914 707162
rect 159294 700718 159326 700954
rect 159562 700718 159646 700954
rect 159882 700718 159914 700954
rect 159294 700634 159914 700718
rect 159294 700398 159326 700634
rect 159562 700398 159646 700634
rect 159882 700398 159914 700634
rect 159294 664954 159914 700398
rect 159294 664718 159326 664954
rect 159562 664718 159646 664954
rect 159882 664718 159914 664954
rect 159294 664634 159914 664718
rect 159294 664398 159326 664634
rect 159562 664398 159646 664634
rect 159882 664398 159914 664634
rect 159294 628954 159914 664398
rect 159294 628718 159326 628954
rect 159562 628718 159646 628954
rect 159882 628718 159914 628954
rect 159294 628634 159914 628718
rect 159294 628398 159326 628634
rect 159562 628398 159646 628634
rect 159882 628398 159914 628634
rect 159294 592954 159914 628398
rect 159294 592718 159326 592954
rect 159562 592718 159646 592954
rect 159882 592718 159914 592954
rect 159294 592634 159914 592718
rect 159294 592398 159326 592634
rect 159562 592398 159646 592634
rect 159882 592398 159914 592634
rect 159294 591292 159914 592398
rect 163794 708678 164414 711590
rect 163794 708442 163826 708678
rect 164062 708442 164146 708678
rect 164382 708442 164414 708678
rect 163794 708358 164414 708442
rect 163794 708122 163826 708358
rect 164062 708122 164146 708358
rect 164382 708122 164414 708358
rect 163794 669454 164414 708122
rect 163794 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 164414 669454
rect 163794 669134 164414 669218
rect 163794 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 164414 669134
rect 163794 633454 164414 668898
rect 163794 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 164414 633454
rect 163794 633134 164414 633218
rect 163794 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 164414 633134
rect 163794 597454 164414 632898
rect 163794 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 164414 597454
rect 163794 597134 164414 597218
rect 163794 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 164414 597134
rect 163794 591292 164414 596898
rect 168294 709638 168914 711590
rect 168294 709402 168326 709638
rect 168562 709402 168646 709638
rect 168882 709402 168914 709638
rect 168294 709318 168914 709402
rect 168294 709082 168326 709318
rect 168562 709082 168646 709318
rect 168882 709082 168914 709318
rect 168294 673954 168914 709082
rect 168294 673718 168326 673954
rect 168562 673718 168646 673954
rect 168882 673718 168914 673954
rect 168294 673634 168914 673718
rect 168294 673398 168326 673634
rect 168562 673398 168646 673634
rect 168882 673398 168914 673634
rect 168294 637954 168914 673398
rect 168294 637718 168326 637954
rect 168562 637718 168646 637954
rect 168882 637718 168914 637954
rect 168294 637634 168914 637718
rect 168294 637398 168326 637634
rect 168562 637398 168646 637634
rect 168882 637398 168914 637634
rect 168294 601954 168914 637398
rect 168294 601718 168326 601954
rect 168562 601718 168646 601954
rect 168882 601718 168914 601954
rect 168294 601634 168914 601718
rect 168294 601398 168326 601634
rect 168562 601398 168646 601634
rect 168882 601398 168914 601634
rect 168294 591292 168914 601398
rect 172794 710598 173414 711590
rect 172794 710362 172826 710598
rect 173062 710362 173146 710598
rect 173382 710362 173414 710598
rect 172794 710278 173414 710362
rect 172794 710042 172826 710278
rect 173062 710042 173146 710278
rect 173382 710042 173414 710278
rect 172794 678454 173414 710042
rect 172794 678218 172826 678454
rect 173062 678218 173146 678454
rect 173382 678218 173414 678454
rect 172794 678134 173414 678218
rect 172794 677898 172826 678134
rect 173062 677898 173146 678134
rect 173382 677898 173414 678134
rect 172794 642454 173414 677898
rect 172794 642218 172826 642454
rect 173062 642218 173146 642454
rect 173382 642218 173414 642454
rect 172794 642134 173414 642218
rect 172794 641898 172826 642134
rect 173062 641898 173146 642134
rect 173382 641898 173414 642134
rect 172794 606454 173414 641898
rect 172794 606218 172826 606454
rect 173062 606218 173146 606454
rect 173382 606218 173414 606454
rect 172794 606134 173414 606218
rect 172794 605898 172826 606134
rect 173062 605898 173146 606134
rect 173382 605898 173414 606134
rect 172794 591292 173414 605898
rect 177294 711558 177914 711590
rect 177294 711322 177326 711558
rect 177562 711322 177646 711558
rect 177882 711322 177914 711558
rect 177294 711238 177914 711322
rect 177294 711002 177326 711238
rect 177562 711002 177646 711238
rect 177882 711002 177914 711238
rect 177294 682954 177914 711002
rect 177294 682718 177326 682954
rect 177562 682718 177646 682954
rect 177882 682718 177914 682954
rect 177294 682634 177914 682718
rect 177294 682398 177326 682634
rect 177562 682398 177646 682634
rect 177882 682398 177914 682634
rect 177294 646954 177914 682398
rect 177294 646718 177326 646954
rect 177562 646718 177646 646954
rect 177882 646718 177914 646954
rect 177294 646634 177914 646718
rect 177294 646398 177326 646634
rect 177562 646398 177646 646634
rect 177882 646398 177914 646634
rect 177294 610954 177914 646398
rect 177294 610718 177326 610954
rect 177562 610718 177646 610954
rect 177882 610718 177914 610954
rect 177294 610634 177914 610718
rect 177294 610398 177326 610634
rect 177562 610398 177646 610634
rect 177882 610398 177914 610634
rect 177294 591292 177914 610398
rect 181794 704838 182414 711590
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 687454 182414 704282
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 651454 182414 686898
rect 181794 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 182414 651454
rect 181794 651134 182414 651218
rect 181794 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 182414 651134
rect 181794 615454 182414 650898
rect 181794 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 182414 615454
rect 181794 615134 182414 615218
rect 181794 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 182414 615134
rect 181794 591292 182414 614898
rect 186294 705798 186914 711590
rect 186294 705562 186326 705798
rect 186562 705562 186646 705798
rect 186882 705562 186914 705798
rect 186294 705478 186914 705562
rect 186294 705242 186326 705478
rect 186562 705242 186646 705478
rect 186882 705242 186914 705478
rect 186294 691954 186914 705242
rect 186294 691718 186326 691954
rect 186562 691718 186646 691954
rect 186882 691718 186914 691954
rect 186294 691634 186914 691718
rect 186294 691398 186326 691634
rect 186562 691398 186646 691634
rect 186882 691398 186914 691634
rect 186294 655954 186914 691398
rect 186294 655718 186326 655954
rect 186562 655718 186646 655954
rect 186882 655718 186914 655954
rect 186294 655634 186914 655718
rect 186294 655398 186326 655634
rect 186562 655398 186646 655634
rect 186882 655398 186914 655634
rect 186294 619954 186914 655398
rect 186294 619718 186326 619954
rect 186562 619718 186646 619954
rect 186882 619718 186914 619954
rect 186294 619634 186914 619718
rect 186294 619398 186326 619634
rect 186562 619398 186646 619634
rect 186882 619398 186914 619634
rect 186294 591292 186914 619398
rect 190794 706758 191414 711590
rect 190794 706522 190826 706758
rect 191062 706522 191146 706758
rect 191382 706522 191414 706758
rect 190794 706438 191414 706522
rect 190794 706202 190826 706438
rect 191062 706202 191146 706438
rect 191382 706202 191414 706438
rect 190794 696454 191414 706202
rect 190794 696218 190826 696454
rect 191062 696218 191146 696454
rect 191382 696218 191414 696454
rect 190794 696134 191414 696218
rect 190794 695898 190826 696134
rect 191062 695898 191146 696134
rect 191382 695898 191414 696134
rect 190794 660454 191414 695898
rect 190794 660218 190826 660454
rect 191062 660218 191146 660454
rect 191382 660218 191414 660454
rect 190794 660134 191414 660218
rect 190794 659898 190826 660134
rect 191062 659898 191146 660134
rect 191382 659898 191414 660134
rect 190794 624454 191414 659898
rect 190794 624218 190826 624454
rect 191062 624218 191146 624454
rect 191382 624218 191414 624454
rect 190794 624134 191414 624218
rect 190794 623898 190826 624134
rect 191062 623898 191146 624134
rect 191382 623898 191414 624134
rect 190794 591292 191414 623898
rect 195294 707718 195914 711590
rect 195294 707482 195326 707718
rect 195562 707482 195646 707718
rect 195882 707482 195914 707718
rect 195294 707398 195914 707482
rect 195294 707162 195326 707398
rect 195562 707162 195646 707398
rect 195882 707162 195914 707398
rect 195294 700954 195914 707162
rect 195294 700718 195326 700954
rect 195562 700718 195646 700954
rect 195882 700718 195914 700954
rect 195294 700634 195914 700718
rect 195294 700398 195326 700634
rect 195562 700398 195646 700634
rect 195882 700398 195914 700634
rect 195294 664954 195914 700398
rect 195294 664718 195326 664954
rect 195562 664718 195646 664954
rect 195882 664718 195914 664954
rect 195294 664634 195914 664718
rect 195294 664398 195326 664634
rect 195562 664398 195646 664634
rect 195882 664398 195914 664634
rect 195294 628954 195914 664398
rect 195294 628718 195326 628954
rect 195562 628718 195646 628954
rect 195882 628718 195914 628954
rect 195294 628634 195914 628718
rect 195294 628398 195326 628634
rect 195562 628398 195646 628634
rect 195882 628398 195914 628634
rect 195294 592954 195914 628398
rect 195294 592718 195326 592954
rect 195562 592718 195646 592954
rect 195882 592718 195914 592954
rect 195294 592634 195914 592718
rect 195294 592398 195326 592634
rect 195562 592398 195646 592634
rect 195882 592398 195914 592634
rect 100272 583954 100620 583986
rect 100272 583718 100328 583954
rect 100564 583718 100620 583954
rect 100272 583634 100620 583718
rect 100272 583398 100328 583634
rect 100564 583398 100620 583634
rect 100272 583366 100620 583398
rect 190440 583954 190788 583986
rect 190440 583718 190496 583954
rect 190732 583718 190788 583954
rect 190440 583634 190788 583718
rect 190440 583398 190496 583634
rect 190732 583398 190788 583634
rect 190440 583366 190788 583398
rect 100952 579454 101300 579486
rect 100952 579218 101008 579454
rect 101244 579218 101300 579454
rect 100952 579134 101300 579218
rect 100952 578898 101008 579134
rect 101244 578898 101300 579134
rect 100952 578866 101300 578898
rect 189760 579454 190108 579486
rect 189760 579218 189816 579454
rect 190052 579218 190108 579454
rect 189760 579134 190108 579218
rect 189760 578898 189816 579134
rect 190052 578898 190108 579134
rect 189760 578866 190108 578898
rect 96294 565718 96326 565954
rect 96562 565718 96646 565954
rect 96882 565718 96914 565954
rect 96294 565634 96914 565718
rect 96294 565398 96326 565634
rect 96562 565398 96646 565634
rect 96882 565398 96914 565634
rect 96294 529954 96914 565398
rect 195294 556954 195914 592398
rect 195294 556718 195326 556954
rect 195562 556718 195646 556954
rect 195882 556718 195914 556954
rect 195294 556634 195914 556718
rect 195294 556398 195326 556634
rect 195562 556398 195646 556634
rect 195882 556398 195914 556634
rect 100272 547954 100620 547986
rect 100272 547718 100328 547954
rect 100564 547718 100620 547954
rect 100272 547634 100620 547718
rect 100272 547398 100328 547634
rect 100564 547398 100620 547634
rect 100272 547366 100620 547398
rect 190440 547954 190788 547986
rect 190440 547718 190496 547954
rect 190732 547718 190788 547954
rect 190440 547634 190788 547718
rect 190440 547398 190496 547634
rect 190732 547398 190788 547634
rect 190440 547366 190788 547398
rect 100952 543454 101300 543486
rect 100952 543218 101008 543454
rect 101244 543218 101300 543454
rect 100952 543134 101300 543218
rect 100952 542898 101008 543134
rect 101244 542898 101300 543134
rect 100952 542866 101300 542898
rect 189760 543454 190108 543486
rect 189760 543218 189816 543454
rect 190052 543218 190108 543454
rect 189760 543134 190108 543218
rect 189760 542898 189816 543134
rect 190052 542898 190108 543134
rect 189760 542866 190108 542898
rect 96294 529718 96326 529954
rect 96562 529718 96646 529954
rect 96882 529718 96914 529954
rect 96294 529634 96914 529718
rect 96294 529398 96326 529634
rect 96562 529398 96646 529634
rect 96882 529398 96914 529634
rect 96294 493954 96914 529398
rect 195294 520954 195914 556398
rect 195294 520718 195326 520954
rect 195562 520718 195646 520954
rect 195882 520718 195914 520954
rect 195294 520634 195914 520718
rect 195294 520398 195326 520634
rect 195562 520398 195646 520634
rect 195882 520398 195914 520634
rect 100272 511954 100620 511986
rect 100272 511718 100328 511954
rect 100564 511718 100620 511954
rect 100272 511634 100620 511718
rect 100272 511398 100328 511634
rect 100564 511398 100620 511634
rect 100272 511366 100620 511398
rect 190440 511954 190788 511986
rect 190440 511718 190496 511954
rect 190732 511718 190788 511954
rect 190440 511634 190788 511718
rect 190440 511398 190496 511634
rect 190732 511398 190788 511634
rect 190440 511366 190788 511398
rect 100952 507454 101300 507486
rect 100952 507218 101008 507454
rect 101244 507218 101300 507454
rect 100952 507134 101300 507218
rect 100952 506898 101008 507134
rect 101244 506898 101300 507134
rect 100952 506866 101300 506898
rect 189760 507454 190108 507486
rect 189760 507218 189816 507454
rect 190052 507218 190108 507454
rect 189760 507134 190108 507218
rect 189760 506898 189816 507134
rect 190052 506898 190108 507134
rect 189760 506866 190108 506898
rect 112928 499590 112988 500106
rect 114288 499590 114348 500106
rect 115376 499590 115436 500106
rect 117688 499590 117748 500106
rect 112928 499530 113098 499590
rect 114288 499530 114386 499590
rect 115376 499530 115490 499590
rect 96294 493718 96326 493954
rect 96562 493718 96646 493954
rect 96882 493718 96914 493954
rect 96294 493634 96914 493718
rect 96294 493398 96326 493634
rect 96562 493398 96646 493634
rect 96882 493398 96914 493634
rect 96294 457954 96914 493398
rect 96294 457718 96326 457954
rect 96562 457718 96646 457954
rect 96882 457718 96914 457954
rect 96294 457634 96914 457718
rect 96294 457398 96326 457634
rect 96562 457398 96646 457634
rect 96882 457398 96914 457634
rect 96294 421954 96914 457398
rect 96294 421718 96326 421954
rect 96562 421718 96646 421954
rect 96882 421718 96914 421954
rect 96294 421634 96914 421718
rect 96294 421398 96326 421634
rect 96562 421398 96646 421634
rect 96882 421398 96914 421634
rect 96294 385954 96914 421398
rect 96294 385718 96326 385954
rect 96562 385718 96646 385954
rect 96882 385718 96914 385954
rect 96294 385634 96914 385718
rect 96294 385398 96326 385634
rect 96562 385398 96646 385634
rect 96882 385398 96914 385634
rect 96294 349954 96914 385398
rect 96294 349718 96326 349954
rect 96562 349718 96646 349954
rect 96882 349718 96914 349954
rect 96294 349634 96914 349718
rect 96294 349398 96326 349634
rect 96562 349398 96646 349634
rect 96882 349398 96914 349634
rect 96294 313954 96914 349398
rect 96294 313718 96326 313954
rect 96562 313718 96646 313954
rect 96882 313718 96914 313954
rect 96294 313634 96914 313718
rect 96294 313398 96326 313634
rect 96562 313398 96646 313634
rect 96882 313398 96914 313634
rect 96294 277954 96914 313398
rect 96294 277718 96326 277954
rect 96562 277718 96646 277954
rect 96882 277718 96914 277954
rect 96294 277634 96914 277718
rect 96294 277398 96326 277634
rect 96562 277398 96646 277634
rect 96882 277398 96914 277634
rect 96294 241954 96914 277398
rect 96294 241718 96326 241954
rect 96562 241718 96646 241954
rect 96882 241718 96914 241954
rect 96294 241634 96914 241718
rect 96294 241398 96326 241634
rect 96562 241398 96646 241634
rect 96882 241398 96914 241634
rect 96294 205954 96914 241398
rect 96294 205718 96326 205954
rect 96562 205718 96646 205954
rect 96882 205718 96914 205954
rect 96294 205634 96914 205718
rect 96294 205398 96326 205634
rect 96562 205398 96646 205634
rect 96882 205398 96914 205634
rect 96294 169954 96914 205398
rect 96294 169718 96326 169954
rect 96562 169718 96646 169954
rect 96882 169718 96914 169954
rect 96294 169634 96914 169718
rect 96294 169398 96326 169634
rect 96562 169398 96646 169634
rect 96882 169398 96914 169634
rect 96294 133954 96914 169398
rect 96294 133718 96326 133954
rect 96562 133718 96646 133954
rect 96882 133718 96914 133954
rect 96294 133634 96914 133718
rect 96294 133398 96326 133634
rect 96562 133398 96646 133634
rect 96882 133398 96914 133634
rect 96294 97954 96914 133398
rect 96294 97718 96326 97954
rect 96562 97718 96646 97954
rect 96882 97718 96914 97954
rect 96294 97634 96914 97718
rect 96294 97398 96326 97634
rect 96562 97398 96646 97634
rect 96882 97398 96914 97634
rect 96294 61954 96914 97398
rect 96294 61718 96326 61954
rect 96562 61718 96646 61954
rect 96882 61718 96914 61954
rect 96294 61634 96914 61718
rect 96294 61398 96326 61634
rect 96562 61398 96646 61634
rect 96882 61398 96914 61634
rect 96294 25954 96914 61398
rect 96294 25718 96326 25954
rect 96562 25718 96646 25954
rect 96882 25718 96914 25954
rect 96294 25634 96914 25718
rect 96294 25398 96326 25634
rect 96562 25398 96646 25634
rect 96882 25398 96914 25634
rect 96294 -5146 96914 25398
rect 96294 -5382 96326 -5146
rect 96562 -5382 96646 -5146
rect 96882 -5382 96914 -5146
rect 96294 -5466 96914 -5382
rect 96294 -5702 96326 -5466
rect 96562 -5702 96646 -5466
rect 96882 -5702 96914 -5466
rect 96294 -7654 96914 -5702
rect 100794 462454 101414 498000
rect 100794 462218 100826 462454
rect 101062 462218 101146 462454
rect 101382 462218 101414 462454
rect 100794 462134 101414 462218
rect 100794 461898 100826 462134
rect 101062 461898 101146 462134
rect 101382 461898 101414 462134
rect 100794 426454 101414 461898
rect 100794 426218 100826 426454
rect 101062 426218 101146 426454
rect 101382 426218 101414 426454
rect 100794 426134 101414 426218
rect 100794 425898 100826 426134
rect 101062 425898 101146 426134
rect 101382 425898 101414 426134
rect 100794 390454 101414 425898
rect 100794 390218 100826 390454
rect 101062 390218 101146 390454
rect 101382 390218 101414 390454
rect 100794 390134 101414 390218
rect 100794 389898 100826 390134
rect 101062 389898 101146 390134
rect 101382 389898 101414 390134
rect 100794 354454 101414 389898
rect 100794 354218 100826 354454
rect 101062 354218 101146 354454
rect 101382 354218 101414 354454
rect 100794 354134 101414 354218
rect 100794 353898 100826 354134
rect 101062 353898 101146 354134
rect 101382 353898 101414 354134
rect 100794 318454 101414 353898
rect 100794 318218 100826 318454
rect 101062 318218 101146 318454
rect 101382 318218 101414 318454
rect 100794 318134 101414 318218
rect 100794 317898 100826 318134
rect 101062 317898 101146 318134
rect 101382 317898 101414 318134
rect 100794 282454 101414 317898
rect 100794 282218 100826 282454
rect 101062 282218 101146 282454
rect 101382 282218 101414 282454
rect 100794 282134 101414 282218
rect 100794 281898 100826 282134
rect 101062 281898 101146 282134
rect 101382 281898 101414 282134
rect 100794 246454 101414 281898
rect 100794 246218 100826 246454
rect 101062 246218 101146 246454
rect 101382 246218 101414 246454
rect 100794 246134 101414 246218
rect 100794 245898 100826 246134
rect 101062 245898 101146 246134
rect 101382 245898 101414 246134
rect 100794 210454 101414 245898
rect 100794 210218 100826 210454
rect 101062 210218 101146 210454
rect 101382 210218 101414 210454
rect 100794 210134 101414 210218
rect 100794 209898 100826 210134
rect 101062 209898 101146 210134
rect 101382 209898 101414 210134
rect 100794 174454 101414 209898
rect 100794 174218 100826 174454
rect 101062 174218 101146 174454
rect 101382 174218 101414 174454
rect 100794 174134 101414 174218
rect 100794 173898 100826 174134
rect 101062 173898 101146 174134
rect 101382 173898 101414 174134
rect 100794 138454 101414 173898
rect 100794 138218 100826 138454
rect 101062 138218 101146 138454
rect 101382 138218 101414 138454
rect 100794 138134 101414 138218
rect 100794 137898 100826 138134
rect 101062 137898 101146 138134
rect 101382 137898 101414 138134
rect 100794 102454 101414 137898
rect 100794 102218 100826 102454
rect 101062 102218 101146 102454
rect 101382 102218 101414 102454
rect 100794 102134 101414 102218
rect 100794 101898 100826 102134
rect 101062 101898 101146 102134
rect 101382 101898 101414 102134
rect 100794 66454 101414 101898
rect 100794 66218 100826 66454
rect 101062 66218 101146 66454
rect 101382 66218 101414 66454
rect 100794 66134 101414 66218
rect 100794 65898 100826 66134
rect 101062 65898 101146 66134
rect 101382 65898 101414 66134
rect 100794 30454 101414 65898
rect 100794 30218 100826 30454
rect 101062 30218 101146 30454
rect 101382 30218 101414 30454
rect 100794 30134 101414 30218
rect 100794 29898 100826 30134
rect 101062 29898 101146 30134
rect 101382 29898 101414 30134
rect 100794 -6106 101414 29898
rect 100794 -6342 100826 -6106
rect 101062 -6342 101146 -6106
rect 101382 -6342 101414 -6106
rect 100794 -6426 101414 -6342
rect 100794 -6662 100826 -6426
rect 101062 -6662 101146 -6426
rect 101382 -6662 101414 -6426
rect 100794 -7654 101414 -6662
rect 105294 466954 105914 498000
rect 105294 466718 105326 466954
rect 105562 466718 105646 466954
rect 105882 466718 105914 466954
rect 105294 466634 105914 466718
rect 105294 466398 105326 466634
rect 105562 466398 105646 466634
rect 105882 466398 105914 466634
rect 105294 430954 105914 466398
rect 105294 430718 105326 430954
rect 105562 430718 105646 430954
rect 105882 430718 105914 430954
rect 105294 430634 105914 430718
rect 105294 430398 105326 430634
rect 105562 430398 105646 430634
rect 105882 430398 105914 430634
rect 105294 394954 105914 430398
rect 105294 394718 105326 394954
rect 105562 394718 105646 394954
rect 105882 394718 105914 394954
rect 105294 394634 105914 394718
rect 105294 394398 105326 394634
rect 105562 394398 105646 394634
rect 105882 394398 105914 394634
rect 105294 358954 105914 394398
rect 105294 358718 105326 358954
rect 105562 358718 105646 358954
rect 105882 358718 105914 358954
rect 105294 358634 105914 358718
rect 105294 358398 105326 358634
rect 105562 358398 105646 358634
rect 105882 358398 105914 358634
rect 105294 322954 105914 358398
rect 105294 322718 105326 322954
rect 105562 322718 105646 322954
rect 105882 322718 105914 322954
rect 105294 322634 105914 322718
rect 105294 322398 105326 322634
rect 105562 322398 105646 322634
rect 105882 322398 105914 322634
rect 105294 286954 105914 322398
rect 105294 286718 105326 286954
rect 105562 286718 105646 286954
rect 105882 286718 105914 286954
rect 105294 286634 105914 286718
rect 105294 286398 105326 286634
rect 105562 286398 105646 286634
rect 105882 286398 105914 286634
rect 105294 250954 105914 286398
rect 105294 250718 105326 250954
rect 105562 250718 105646 250954
rect 105882 250718 105914 250954
rect 105294 250634 105914 250718
rect 105294 250398 105326 250634
rect 105562 250398 105646 250634
rect 105882 250398 105914 250634
rect 105294 214954 105914 250398
rect 105294 214718 105326 214954
rect 105562 214718 105646 214954
rect 105882 214718 105914 214954
rect 105294 214634 105914 214718
rect 105294 214398 105326 214634
rect 105562 214398 105646 214634
rect 105882 214398 105914 214634
rect 105294 178954 105914 214398
rect 105294 178718 105326 178954
rect 105562 178718 105646 178954
rect 105882 178718 105914 178954
rect 105294 178634 105914 178718
rect 105294 178398 105326 178634
rect 105562 178398 105646 178634
rect 105882 178398 105914 178634
rect 105294 142954 105914 178398
rect 105294 142718 105326 142954
rect 105562 142718 105646 142954
rect 105882 142718 105914 142954
rect 105294 142634 105914 142718
rect 105294 142398 105326 142634
rect 105562 142398 105646 142634
rect 105882 142398 105914 142634
rect 105294 106954 105914 142398
rect 105294 106718 105326 106954
rect 105562 106718 105646 106954
rect 105882 106718 105914 106954
rect 105294 106634 105914 106718
rect 105294 106398 105326 106634
rect 105562 106398 105646 106634
rect 105882 106398 105914 106634
rect 105294 70954 105914 106398
rect 105294 70718 105326 70954
rect 105562 70718 105646 70954
rect 105882 70718 105914 70954
rect 105294 70634 105914 70718
rect 105294 70398 105326 70634
rect 105562 70398 105646 70634
rect 105882 70398 105914 70634
rect 105294 34954 105914 70398
rect 105294 34718 105326 34954
rect 105562 34718 105646 34954
rect 105882 34718 105914 34954
rect 105294 34634 105914 34718
rect 105294 34398 105326 34634
rect 105562 34398 105646 34634
rect 105882 34398 105914 34634
rect 105294 -7066 105914 34398
rect 105294 -7302 105326 -7066
rect 105562 -7302 105646 -7066
rect 105882 -7302 105914 -7066
rect 105294 -7386 105914 -7302
rect 105294 -7622 105326 -7386
rect 105562 -7622 105646 -7386
rect 105882 -7622 105914 -7386
rect 105294 -7654 105914 -7622
rect 109794 471454 110414 498000
rect 113038 496909 113098 499530
rect 114326 498269 114386 499530
rect 114323 498268 114389 498269
rect 114323 498204 114324 498268
rect 114388 498204 114389 498268
rect 114323 498203 114389 498204
rect 113035 496908 113101 496909
rect 113035 496844 113036 496908
rect 113100 496844 113101 496908
rect 113035 496843 113101 496844
rect 109794 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 110414 471454
rect 109794 471134 110414 471218
rect 109794 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 110414 471134
rect 109794 435454 110414 470898
rect 109794 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 110414 435454
rect 109794 435134 110414 435218
rect 109794 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 110414 435134
rect 109794 399454 110414 434898
rect 109794 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 110414 399454
rect 109794 399134 110414 399218
rect 109794 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 110414 399134
rect 109794 363454 110414 398898
rect 109794 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 110414 363454
rect 109794 363134 110414 363218
rect 109794 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 110414 363134
rect 109794 327454 110414 362898
rect 109794 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 110414 327454
rect 109794 327134 110414 327218
rect 109794 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 110414 327134
rect 109794 291454 110414 326898
rect 109794 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 110414 291454
rect 109794 291134 110414 291218
rect 109794 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 110414 291134
rect 109794 255454 110414 290898
rect 109794 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 110414 255454
rect 109794 255134 110414 255218
rect 109794 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 110414 255134
rect 109794 219454 110414 254898
rect 109794 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 110414 219454
rect 109794 219134 110414 219218
rect 109794 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 110414 219134
rect 109794 183454 110414 218898
rect 109794 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 110414 183454
rect 109794 183134 110414 183218
rect 109794 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 110414 183134
rect 109794 147454 110414 182898
rect 109794 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 110414 147454
rect 109794 147134 110414 147218
rect 109794 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 110414 147134
rect 109794 111454 110414 146898
rect 109794 111218 109826 111454
rect 110062 111218 110146 111454
rect 110382 111218 110414 111454
rect 109794 111134 110414 111218
rect 109794 110898 109826 111134
rect 110062 110898 110146 111134
rect 110382 110898 110414 111134
rect 109794 75454 110414 110898
rect 109794 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 110414 75454
rect 109794 75134 110414 75218
rect 109794 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 110414 75134
rect 109794 39454 110414 74898
rect 109794 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 110414 39454
rect 109794 39134 110414 39218
rect 109794 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 110414 39134
rect 109794 3454 110414 38898
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -7654 110414 -902
rect 114294 475954 114914 498000
rect 115430 496909 115490 499530
rect 117638 499530 117748 499590
rect 118912 499590 118972 500106
rect 120000 499590 120060 500106
rect 121088 499590 121148 500106
rect 122312 499590 122372 500106
rect 123400 499590 123460 500106
rect 118912 499530 118986 499590
rect 120000 499530 120090 499590
rect 121088 499530 121194 499590
rect 122312 499530 122482 499590
rect 117638 496909 117698 499530
rect 118926 498269 118986 499530
rect 118923 498268 118989 498269
rect 118923 498204 118924 498268
rect 118988 498204 118989 498268
rect 118923 498203 118989 498204
rect 115427 496908 115493 496909
rect 115427 496844 115428 496908
rect 115492 496844 115493 496908
rect 115427 496843 115493 496844
rect 117635 496908 117701 496909
rect 117635 496844 117636 496908
rect 117700 496844 117701 496908
rect 117635 496843 117701 496844
rect 114294 475718 114326 475954
rect 114562 475718 114646 475954
rect 114882 475718 114914 475954
rect 114294 475634 114914 475718
rect 114294 475398 114326 475634
rect 114562 475398 114646 475634
rect 114882 475398 114914 475634
rect 114294 439954 114914 475398
rect 114294 439718 114326 439954
rect 114562 439718 114646 439954
rect 114882 439718 114914 439954
rect 114294 439634 114914 439718
rect 114294 439398 114326 439634
rect 114562 439398 114646 439634
rect 114882 439398 114914 439634
rect 114294 403954 114914 439398
rect 114294 403718 114326 403954
rect 114562 403718 114646 403954
rect 114882 403718 114914 403954
rect 114294 403634 114914 403718
rect 114294 403398 114326 403634
rect 114562 403398 114646 403634
rect 114882 403398 114914 403634
rect 114294 367954 114914 403398
rect 114294 367718 114326 367954
rect 114562 367718 114646 367954
rect 114882 367718 114914 367954
rect 114294 367634 114914 367718
rect 114294 367398 114326 367634
rect 114562 367398 114646 367634
rect 114882 367398 114914 367634
rect 114294 331954 114914 367398
rect 114294 331718 114326 331954
rect 114562 331718 114646 331954
rect 114882 331718 114914 331954
rect 114294 331634 114914 331718
rect 114294 331398 114326 331634
rect 114562 331398 114646 331634
rect 114882 331398 114914 331634
rect 114294 295954 114914 331398
rect 114294 295718 114326 295954
rect 114562 295718 114646 295954
rect 114882 295718 114914 295954
rect 114294 295634 114914 295718
rect 114294 295398 114326 295634
rect 114562 295398 114646 295634
rect 114882 295398 114914 295634
rect 114294 259954 114914 295398
rect 114294 259718 114326 259954
rect 114562 259718 114646 259954
rect 114882 259718 114914 259954
rect 114294 259634 114914 259718
rect 114294 259398 114326 259634
rect 114562 259398 114646 259634
rect 114882 259398 114914 259634
rect 114294 223954 114914 259398
rect 114294 223718 114326 223954
rect 114562 223718 114646 223954
rect 114882 223718 114914 223954
rect 114294 223634 114914 223718
rect 114294 223398 114326 223634
rect 114562 223398 114646 223634
rect 114882 223398 114914 223634
rect 114294 187954 114914 223398
rect 114294 187718 114326 187954
rect 114562 187718 114646 187954
rect 114882 187718 114914 187954
rect 114294 187634 114914 187718
rect 114294 187398 114326 187634
rect 114562 187398 114646 187634
rect 114882 187398 114914 187634
rect 114294 151954 114914 187398
rect 114294 151718 114326 151954
rect 114562 151718 114646 151954
rect 114882 151718 114914 151954
rect 114294 151634 114914 151718
rect 114294 151398 114326 151634
rect 114562 151398 114646 151634
rect 114882 151398 114914 151634
rect 114294 115954 114914 151398
rect 114294 115718 114326 115954
rect 114562 115718 114646 115954
rect 114882 115718 114914 115954
rect 114294 115634 114914 115718
rect 114294 115398 114326 115634
rect 114562 115398 114646 115634
rect 114882 115398 114914 115634
rect 114294 79954 114914 115398
rect 114294 79718 114326 79954
rect 114562 79718 114646 79954
rect 114882 79718 114914 79954
rect 114294 79634 114914 79718
rect 114294 79398 114326 79634
rect 114562 79398 114646 79634
rect 114882 79398 114914 79634
rect 114294 43954 114914 79398
rect 114294 43718 114326 43954
rect 114562 43718 114646 43954
rect 114882 43718 114914 43954
rect 114294 43634 114914 43718
rect 114294 43398 114326 43634
rect 114562 43398 114646 43634
rect 114882 43398 114914 43634
rect 114294 7954 114914 43398
rect 114294 7718 114326 7954
rect 114562 7718 114646 7954
rect 114882 7718 114914 7954
rect 114294 7634 114914 7718
rect 114294 7398 114326 7634
rect 114562 7398 114646 7634
rect 114882 7398 114914 7634
rect 114294 -1306 114914 7398
rect 114294 -1542 114326 -1306
rect 114562 -1542 114646 -1306
rect 114882 -1542 114914 -1306
rect 114294 -1626 114914 -1542
rect 114294 -1862 114326 -1626
rect 114562 -1862 114646 -1626
rect 114882 -1862 114914 -1626
rect 114294 -7654 114914 -1862
rect 118794 480454 119414 498000
rect 120030 497453 120090 499530
rect 120027 497452 120093 497453
rect 120027 497388 120028 497452
rect 120092 497388 120093 497452
rect 120027 497387 120093 497388
rect 121134 496909 121194 499530
rect 122422 496909 122482 499530
rect 123342 499530 123460 499590
rect 124760 499590 124820 500106
rect 125304 499590 125364 500106
rect 125712 499590 125772 500106
rect 130472 499590 130532 500106
rect 135504 499590 135564 500106
rect 124760 499530 124874 499590
rect 125304 499530 125426 499590
rect 125712 499530 125794 499590
rect 130472 499530 130578 499590
rect 123342 498269 123402 499530
rect 123339 498268 123405 498269
rect 123339 498204 123340 498268
rect 123404 498204 123405 498268
rect 123339 498203 123405 498204
rect 124814 498133 124874 499530
rect 124811 498132 124877 498133
rect 124811 498068 124812 498132
rect 124876 498068 124877 498132
rect 124811 498067 124877 498068
rect 121131 496908 121197 496909
rect 121131 496844 121132 496908
rect 121196 496844 121197 496908
rect 121131 496843 121197 496844
rect 122419 496908 122485 496909
rect 122419 496844 122420 496908
rect 122484 496844 122485 496908
rect 122419 496843 122485 496844
rect 118794 480218 118826 480454
rect 119062 480218 119146 480454
rect 119382 480218 119414 480454
rect 118794 480134 119414 480218
rect 118794 479898 118826 480134
rect 119062 479898 119146 480134
rect 119382 479898 119414 480134
rect 118794 444454 119414 479898
rect 118794 444218 118826 444454
rect 119062 444218 119146 444454
rect 119382 444218 119414 444454
rect 118794 444134 119414 444218
rect 118794 443898 118826 444134
rect 119062 443898 119146 444134
rect 119382 443898 119414 444134
rect 118794 408454 119414 443898
rect 118794 408218 118826 408454
rect 119062 408218 119146 408454
rect 119382 408218 119414 408454
rect 118794 408134 119414 408218
rect 118794 407898 118826 408134
rect 119062 407898 119146 408134
rect 119382 407898 119414 408134
rect 118794 372454 119414 407898
rect 118794 372218 118826 372454
rect 119062 372218 119146 372454
rect 119382 372218 119414 372454
rect 118794 372134 119414 372218
rect 118794 371898 118826 372134
rect 119062 371898 119146 372134
rect 119382 371898 119414 372134
rect 118794 336454 119414 371898
rect 118794 336218 118826 336454
rect 119062 336218 119146 336454
rect 119382 336218 119414 336454
rect 118794 336134 119414 336218
rect 118794 335898 118826 336134
rect 119062 335898 119146 336134
rect 119382 335898 119414 336134
rect 118794 300454 119414 335898
rect 118794 300218 118826 300454
rect 119062 300218 119146 300454
rect 119382 300218 119414 300454
rect 118794 300134 119414 300218
rect 118794 299898 118826 300134
rect 119062 299898 119146 300134
rect 119382 299898 119414 300134
rect 118794 264454 119414 299898
rect 118794 264218 118826 264454
rect 119062 264218 119146 264454
rect 119382 264218 119414 264454
rect 118794 264134 119414 264218
rect 118794 263898 118826 264134
rect 119062 263898 119146 264134
rect 119382 263898 119414 264134
rect 118794 228454 119414 263898
rect 118794 228218 118826 228454
rect 119062 228218 119146 228454
rect 119382 228218 119414 228454
rect 118794 228134 119414 228218
rect 118794 227898 118826 228134
rect 119062 227898 119146 228134
rect 119382 227898 119414 228134
rect 118794 192454 119414 227898
rect 118794 192218 118826 192454
rect 119062 192218 119146 192454
rect 119382 192218 119414 192454
rect 118794 192134 119414 192218
rect 118794 191898 118826 192134
rect 119062 191898 119146 192134
rect 119382 191898 119414 192134
rect 118794 156454 119414 191898
rect 118794 156218 118826 156454
rect 119062 156218 119146 156454
rect 119382 156218 119414 156454
rect 118794 156134 119414 156218
rect 118794 155898 118826 156134
rect 119062 155898 119146 156134
rect 119382 155898 119414 156134
rect 118794 120454 119414 155898
rect 118794 120218 118826 120454
rect 119062 120218 119146 120454
rect 119382 120218 119414 120454
rect 118794 120134 119414 120218
rect 118794 119898 118826 120134
rect 119062 119898 119146 120134
rect 119382 119898 119414 120134
rect 118794 84454 119414 119898
rect 118794 84218 118826 84454
rect 119062 84218 119146 84454
rect 119382 84218 119414 84454
rect 118794 84134 119414 84218
rect 118794 83898 118826 84134
rect 119062 83898 119146 84134
rect 119382 83898 119414 84134
rect 118794 48454 119414 83898
rect 118794 48218 118826 48454
rect 119062 48218 119146 48454
rect 119382 48218 119414 48454
rect 118794 48134 119414 48218
rect 118794 47898 118826 48134
rect 119062 47898 119146 48134
rect 119382 47898 119414 48134
rect 118794 12454 119414 47898
rect 118794 12218 118826 12454
rect 119062 12218 119146 12454
rect 119382 12218 119414 12454
rect 118794 12134 119414 12218
rect 118794 11898 118826 12134
rect 119062 11898 119146 12134
rect 119382 11898 119414 12134
rect 118794 -2266 119414 11898
rect 118794 -2502 118826 -2266
rect 119062 -2502 119146 -2266
rect 119382 -2502 119414 -2266
rect 118794 -2586 119414 -2502
rect 118794 -2822 118826 -2586
rect 119062 -2822 119146 -2586
rect 119382 -2822 119414 -2586
rect 118794 -7654 119414 -2822
rect 123294 484954 123914 498000
rect 125366 496909 125426 499530
rect 125734 498133 125794 499530
rect 125731 498132 125797 498133
rect 125731 498068 125732 498132
rect 125796 498068 125797 498132
rect 125731 498067 125797 498068
rect 125363 496908 125429 496909
rect 125363 496844 125364 496908
rect 125428 496844 125429 496908
rect 125363 496843 125429 496844
rect 123294 484718 123326 484954
rect 123562 484718 123646 484954
rect 123882 484718 123914 484954
rect 123294 484634 123914 484718
rect 123294 484398 123326 484634
rect 123562 484398 123646 484634
rect 123882 484398 123914 484634
rect 123294 448954 123914 484398
rect 123294 448718 123326 448954
rect 123562 448718 123646 448954
rect 123882 448718 123914 448954
rect 123294 448634 123914 448718
rect 123294 448398 123326 448634
rect 123562 448398 123646 448634
rect 123882 448398 123914 448634
rect 123294 412954 123914 448398
rect 123294 412718 123326 412954
rect 123562 412718 123646 412954
rect 123882 412718 123914 412954
rect 123294 412634 123914 412718
rect 123294 412398 123326 412634
rect 123562 412398 123646 412634
rect 123882 412398 123914 412634
rect 123294 376954 123914 412398
rect 123294 376718 123326 376954
rect 123562 376718 123646 376954
rect 123882 376718 123914 376954
rect 123294 376634 123914 376718
rect 123294 376398 123326 376634
rect 123562 376398 123646 376634
rect 123882 376398 123914 376634
rect 123294 340954 123914 376398
rect 123294 340718 123326 340954
rect 123562 340718 123646 340954
rect 123882 340718 123914 340954
rect 123294 340634 123914 340718
rect 123294 340398 123326 340634
rect 123562 340398 123646 340634
rect 123882 340398 123914 340634
rect 123294 304954 123914 340398
rect 123294 304718 123326 304954
rect 123562 304718 123646 304954
rect 123882 304718 123914 304954
rect 123294 304634 123914 304718
rect 123294 304398 123326 304634
rect 123562 304398 123646 304634
rect 123882 304398 123914 304634
rect 123294 268954 123914 304398
rect 123294 268718 123326 268954
rect 123562 268718 123646 268954
rect 123882 268718 123914 268954
rect 123294 268634 123914 268718
rect 123294 268398 123326 268634
rect 123562 268398 123646 268634
rect 123882 268398 123914 268634
rect 123294 232954 123914 268398
rect 123294 232718 123326 232954
rect 123562 232718 123646 232954
rect 123882 232718 123914 232954
rect 123294 232634 123914 232718
rect 123294 232398 123326 232634
rect 123562 232398 123646 232634
rect 123882 232398 123914 232634
rect 123294 196954 123914 232398
rect 123294 196718 123326 196954
rect 123562 196718 123646 196954
rect 123882 196718 123914 196954
rect 123294 196634 123914 196718
rect 123294 196398 123326 196634
rect 123562 196398 123646 196634
rect 123882 196398 123914 196634
rect 123294 160954 123914 196398
rect 123294 160718 123326 160954
rect 123562 160718 123646 160954
rect 123882 160718 123914 160954
rect 123294 160634 123914 160718
rect 123294 160398 123326 160634
rect 123562 160398 123646 160634
rect 123882 160398 123914 160634
rect 123294 124954 123914 160398
rect 123294 124718 123326 124954
rect 123562 124718 123646 124954
rect 123882 124718 123914 124954
rect 123294 124634 123914 124718
rect 123294 124398 123326 124634
rect 123562 124398 123646 124634
rect 123882 124398 123914 124634
rect 123294 88954 123914 124398
rect 123294 88718 123326 88954
rect 123562 88718 123646 88954
rect 123882 88718 123914 88954
rect 123294 88634 123914 88718
rect 123294 88398 123326 88634
rect 123562 88398 123646 88634
rect 123882 88398 123914 88634
rect 123294 52954 123914 88398
rect 123294 52718 123326 52954
rect 123562 52718 123646 52954
rect 123882 52718 123914 52954
rect 123294 52634 123914 52718
rect 123294 52398 123326 52634
rect 123562 52398 123646 52634
rect 123882 52398 123914 52634
rect 123294 16954 123914 52398
rect 123294 16718 123326 16954
rect 123562 16718 123646 16954
rect 123882 16718 123914 16954
rect 123294 16634 123914 16718
rect 123294 16398 123326 16634
rect 123562 16398 123646 16634
rect 123882 16398 123914 16634
rect 123294 -3226 123914 16398
rect 123294 -3462 123326 -3226
rect 123562 -3462 123646 -3226
rect 123882 -3462 123914 -3226
rect 123294 -3546 123914 -3462
rect 123294 -3782 123326 -3546
rect 123562 -3782 123646 -3546
rect 123882 -3782 123914 -3546
rect 123294 -7654 123914 -3782
rect 127794 489454 128414 498000
rect 130518 496909 130578 499530
rect 135486 499530 135564 499590
rect 140536 499590 140596 500106
rect 145568 499590 145628 500106
rect 150464 499590 150524 500106
rect 155496 499590 155556 500106
rect 160528 499590 160588 500106
rect 140536 499530 140698 499590
rect 145568 499530 145666 499590
rect 150464 499530 150634 499590
rect 155496 499530 155602 499590
rect 130515 496908 130581 496909
rect 130515 496844 130516 496908
rect 130580 496844 130581 496908
rect 130515 496843 130581 496844
rect 127794 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 128414 489454
rect 127794 489134 128414 489218
rect 127794 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 128414 489134
rect 127794 453454 128414 488898
rect 127794 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 128414 453454
rect 127794 453134 128414 453218
rect 127794 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 128414 453134
rect 127794 417454 128414 452898
rect 127794 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 128414 417454
rect 127794 417134 128414 417218
rect 127794 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 128414 417134
rect 127794 381454 128414 416898
rect 127794 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 128414 381454
rect 127794 381134 128414 381218
rect 127794 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 128414 381134
rect 127794 345454 128414 380898
rect 127794 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 128414 345454
rect 127794 345134 128414 345218
rect 127794 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 128414 345134
rect 127794 309454 128414 344898
rect 127794 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 128414 309454
rect 127794 309134 128414 309218
rect 127794 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 128414 309134
rect 127794 273454 128414 308898
rect 127794 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 128414 273454
rect 127794 273134 128414 273218
rect 127794 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 128414 273134
rect 127794 237454 128414 272898
rect 127794 237218 127826 237454
rect 128062 237218 128146 237454
rect 128382 237218 128414 237454
rect 127794 237134 128414 237218
rect 127794 236898 127826 237134
rect 128062 236898 128146 237134
rect 128382 236898 128414 237134
rect 127794 201454 128414 236898
rect 127794 201218 127826 201454
rect 128062 201218 128146 201454
rect 128382 201218 128414 201454
rect 127794 201134 128414 201218
rect 127794 200898 127826 201134
rect 128062 200898 128146 201134
rect 128382 200898 128414 201134
rect 127794 165454 128414 200898
rect 127794 165218 127826 165454
rect 128062 165218 128146 165454
rect 128382 165218 128414 165454
rect 127794 165134 128414 165218
rect 127794 164898 127826 165134
rect 128062 164898 128146 165134
rect 128382 164898 128414 165134
rect 127794 129454 128414 164898
rect 127794 129218 127826 129454
rect 128062 129218 128146 129454
rect 128382 129218 128414 129454
rect 127794 129134 128414 129218
rect 127794 128898 127826 129134
rect 128062 128898 128146 129134
rect 128382 128898 128414 129134
rect 127794 93454 128414 128898
rect 127794 93218 127826 93454
rect 128062 93218 128146 93454
rect 128382 93218 128414 93454
rect 127794 93134 128414 93218
rect 127794 92898 127826 93134
rect 128062 92898 128146 93134
rect 128382 92898 128414 93134
rect 127794 57454 128414 92898
rect 127794 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 128414 57454
rect 127794 57134 128414 57218
rect 127794 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 128414 57134
rect 127794 21454 128414 56898
rect 127794 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 128414 21454
rect 127794 21134 128414 21218
rect 127794 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 128414 21134
rect 127794 -4186 128414 20898
rect 127794 -4422 127826 -4186
rect 128062 -4422 128146 -4186
rect 128382 -4422 128414 -4186
rect 127794 -4506 128414 -4422
rect 127794 -4742 127826 -4506
rect 128062 -4742 128146 -4506
rect 128382 -4742 128414 -4506
rect 127794 -7654 128414 -4742
rect 132294 493954 132914 498000
rect 135486 496909 135546 499530
rect 135483 496908 135549 496909
rect 135483 496844 135484 496908
rect 135548 496844 135549 496908
rect 135483 496843 135549 496844
rect 132294 493718 132326 493954
rect 132562 493718 132646 493954
rect 132882 493718 132914 493954
rect 132294 493634 132914 493718
rect 132294 493398 132326 493634
rect 132562 493398 132646 493634
rect 132882 493398 132914 493634
rect 132294 457954 132914 493398
rect 132294 457718 132326 457954
rect 132562 457718 132646 457954
rect 132882 457718 132914 457954
rect 132294 457634 132914 457718
rect 132294 457398 132326 457634
rect 132562 457398 132646 457634
rect 132882 457398 132914 457634
rect 132294 421954 132914 457398
rect 132294 421718 132326 421954
rect 132562 421718 132646 421954
rect 132882 421718 132914 421954
rect 132294 421634 132914 421718
rect 132294 421398 132326 421634
rect 132562 421398 132646 421634
rect 132882 421398 132914 421634
rect 132294 385954 132914 421398
rect 132294 385718 132326 385954
rect 132562 385718 132646 385954
rect 132882 385718 132914 385954
rect 132294 385634 132914 385718
rect 132294 385398 132326 385634
rect 132562 385398 132646 385634
rect 132882 385398 132914 385634
rect 132294 349954 132914 385398
rect 132294 349718 132326 349954
rect 132562 349718 132646 349954
rect 132882 349718 132914 349954
rect 132294 349634 132914 349718
rect 132294 349398 132326 349634
rect 132562 349398 132646 349634
rect 132882 349398 132914 349634
rect 132294 313954 132914 349398
rect 132294 313718 132326 313954
rect 132562 313718 132646 313954
rect 132882 313718 132914 313954
rect 132294 313634 132914 313718
rect 132294 313398 132326 313634
rect 132562 313398 132646 313634
rect 132882 313398 132914 313634
rect 132294 277954 132914 313398
rect 132294 277718 132326 277954
rect 132562 277718 132646 277954
rect 132882 277718 132914 277954
rect 132294 277634 132914 277718
rect 132294 277398 132326 277634
rect 132562 277398 132646 277634
rect 132882 277398 132914 277634
rect 132294 241954 132914 277398
rect 132294 241718 132326 241954
rect 132562 241718 132646 241954
rect 132882 241718 132914 241954
rect 132294 241634 132914 241718
rect 132294 241398 132326 241634
rect 132562 241398 132646 241634
rect 132882 241398 132914 241634
rect 132294 205954 132914 241398
rect 132294 205718 132326 205954
rect 132562 205718 132646 205954
rect 132882 205718 132914 205954
rect 132294 205634 132914 205718
rect 132294 205398 132326 205634
rect 132562 205398 132646 205634
rect 132882 205398 132914 205634
rect 132294 169954 132914 205398
rect 132294 169718 132326 169954
rect 132562 169718 132646 169954
rect 132882 169718 132914 169954
rect 132294 169634 132914 169718
rect 132294 169398 132326 169634
rect 132562 169398 132646 169634
rect 132882 169398 132914 169634
rect 132294 133954 132914 169398
rect 132294 133718 132326 133954
rect 132562 133718 132646 133954
rect 132882 133718 132914 133954
rect 132294 133634 132914 133718
rect 132294 133398 132326 133634
rect 132562 133398 132646 133634
rect 132882 133398 132914 133634
rect 132294 97954 132914 133398
rect 132294 97718 132326 97954
rect 132562 97718 132646 97954
rect 132882 97718 132914 97954
rect 132294 97634 132914 97718
rect 132294 97398 132326 97634
rect 132562 97398 132646 97634
rect 132882 97398 132914 97634
rect 132294 61954 132914 97398
rect 132294 61718 132326 61954
rect 132562 61718 132646 61954
rect 132882 61718 132914 61954
rect 132294 61634 132914 61718
rect 132294 61398 132326 61634
rect 132562 61398 132646 61634
rect 132882 61398 132914 61634
rect 132294 25954 132914 61398
rect 132294 25718 132326 25954
rect 132562 25718 132646 25954
rect 132882 25718 132914 25954
rect 132294 25634 132914 25718
rect 132294 25398 132326 25634
rect 132562 25398 132646 25634
rect 132882 25398 132914 25634
rect 132294 -5146 132914 25398
rect 132294 -5382 132326 -5146
rect 132562 -5382 132646 -5146
rect 132882 -5382 132914 -5146
rect 132294 -5466 132914 -5382
rect 132294 -5702 132326 -5466
rect 132562 -5702 132646 -5466
rect 132882 -5702 132914 -5466
rect 132294 -7654 132914 -5702
rect 136794 462454 137414 498000
rect 140638 496909 140698 499530
rect 140635 496908 140701 496909
rect 140635 496844 140636 496908
rect 140700 496844 140701 496908
rect 140635 496843 140701 496844
rect 136794 462218 136826 462454
rect 137062 462218 137146 462454
rect 137382 462218 137414 462454
rect 136794 462134 137414 462218
rect 136794 461898 136826 462134
rect 137062 461898 137146 462134
rect 137382 461898 137414 462134
rect 136794 426454 137414 461898
rect 136794 426218 136826 426454
rect 137062 426218 137146 426454
rect 137382 426218 137414 426454
rect 136794 426134 137414 426218
rect 136794 425898 136826 426134
rect 137062 425898 137146 426134
rect 137382 425898 137414 426134
rect 136794 390454 137414 425898
rect 136794 390218 136826 390454
rect 137062 390218 137146 390454
rect 137382 390218 137414 390454
rect 136794 390134 137414 390218
rect 136794 389898 136826 390134
rect 137062 389898 137146 390134
rect 137382 389898 137414 390134
rect 136794 354454 137414 389898
rect 136794 354218 136826 354454
rect 137062 354218 137146 354454
rect 137382 354218 137414 354454
rect 136794 354134 137414 354218
rect 136794 353898 136826 354134
rect 137062 353898 137146 354134
rect 137382 353898 137414 354134
rect 136794 318454 137414 353898
rect 136794 318218 136826 318454
rect 137062 318218 137146 318454
rect 137382 318218 137414 318454
rect 136794 318134 137414 318218
rect 136794 317898 136826 318134
rect 137062 317898 137146 318134
rect 137382 317898 137414 318134
rect 136794 282454 137414 317898
rect 136794 282218 136826 282454
rect 137062 282218 137146 282454
rect 137382 282218 137414 282454
rect 136794 282134 137414 282218
rect 136794 281898 136826 282134
rect 137062 281898 137146 282134
rect 137382 281898 137414 282134
rect 136794 246454 137414 281898
rect 136794 246218 136826 246454
rect 137062 246218 137146 246454
rect 137382 246218 137414 246454
rect 136794 246134 137414 246218
rect 136794 245898 136826 246134
rect 137062 245898 137146 246134
rect 137382 245898 137414 246134
rect 136794 210454 137414 245898
rect 136794 210218 136826 210454
rect 137062 210218 137146 210454
rect 137382 210218 137414 210454
rect 136794 210134 137414 210218
rect 136794 209898 136826 210134
rect 137062 209898 137146 210134
rect 137382 209898 137414 210134
rect 136794 174454 137414 209898
rect 136794 174218 136826 174454
rect 137062 174218 137146 174454
rect 137382 174218 137414 174454
rect 136794 174134 137414 174218
rect 136794 173898 136826 174134
rect 137062 173898 137146 174134
rect 137382 173898 137414 174134
rect 136794 138454 137414 173898
rect 136794 138218 136826 138454
rect 137062 138218 137146 138454
rect 137382 138218 137414 138454
rect 136794 138134 137414 138218
rect 136794 137898 136826 138134
rect 137062 137898 137146 138134
rect 137382 137898 137414 138134
rect 136794 102454 137414 137898
rect 136794 102218 136826 102454
rect 137062 102218 137146 102454
rect 137382 102218 137414 102454
rect 136794 102134 137414 102218
rect 136794 101898 136826 102134
rect 137062 101898 137146 102134
rect 137382 101898 137414 102134
rect 136794 66454 137414 101898
rect 136794 66218 136826 66454
rect 137062 66218 137146 66454
rect 137382 66218 137414 66454
rect 136794 66134 137414 66218
rect 136794 65898 136826 66134
rect 137062 65898 137146 66134
rect 137382 65898 137414 66134
rect 136794 30454 137414 65898
rect 136794 30218 136826 30454
rect 137062 30218 137146 30454
rect 137382 30218 137414 30454
rect 136794 30134 137414 30218
rect 136794 29898 136826 30134
rect 137062 29898 137146 30134
rect 137382 29898 137414 30134
rect 136794 -6106 137414 29898
rect 136794 -6342 136826 -6106
rect 137062 -6342 137146 -6106
rect 137382 -6342 137414 -6106
rect 136794 -6426 137414 -6342
rect 136794 -6662 136826 -6426
rect 137062 -6662 137146 -6426
rect 137382 -6662 137414 -6426
rect 136794 -7654 137414 -6662
rect 141294 466954 141914 498000
rect 145606 496909 145666 499530
rect 150574 498269 150634 499530
rect 150571 498268 150637 498269
rect 150571 498204 150572 498268
rect 150636 498204 150637 498268
rect 150571 498203 150637 498204
rect 145603 496908 145669 496909
rect 145603 496844 145604 496908
rect 145668 496844 145669 496908
rect 145603 496843 145669 496844
rect 141294 466718 141326 466954
rect 141562 466718 141646 466954
rect 141882 466718 141914 466954
rect 141294 466634 141914 466718
rect 141294 466398 141326 466634
rect 141562 466398 141646 466634
rect 141882 466398 141914 466634
rect 141294 430954 141914 466398
rect 141294 430718 141326 430954
rect 141562 430718 141646 430954
rect 141882 430718 141914 430954
rect 141294 430634 141914 430718
rect 141294 430398 141326 430634
rect 141562 430398 141646 430634
rect 141882 430398 141914 430634
rect 141294 394954 141914 430398
rect 141294 394718 141326 394954
rect 141562 394718 141646 394954
rect 141882 394718 141914 394954
rect 141294 394634 141914 394718
rect 141294 394398 141326 394634
rect 141562 394398 141646 394634
rect 141882 394398 141914 394634
rect 141294 358954 141914 394398
rect 141294 358718 141326 358954
rect 141562 358718 141646 358954
rect 141882 358718 141914 358954
rect 141294 358634 141914 358718
rect 141294 358398 141326 358634
rect 141562 358398 141646 358634
rect 141882 358398 141914 358634
rect 141294 322954 141914 358398
rect 141294 322718 141326 322954
rect 141562 322718 141646 322954
rect 141882 322718 141914 322954
rect 141294 322634 141914 322718
rect 141294 322398 141326 322634
rect 141562 322398 141646 322634
rect 141882 322398 141914 322634
rect 141294 286954 141914 322398
rect 141294 286718 141326 286954
rect 141562 286718 141646 286954
rect 141882 286718 141914 286954
rect 141294 286634 141914 286718
rect 141294 286398 141326 286634
rect 141562 286398 141646 286634
rect 141882 286398 141914 286634
rect 141294 250954 141914 286398
rect 141294 250718 141326 250954
rect 141562 250718 141646 250954
rect 141882 250718 141914 250954
rect 141294 250634 141914 250718
rect 141294 250398 141326 250634
rect 141562 250398 141646 250634
rect 141882 250398 141914 250634
rect 141294 214954 141914 250398
rect 141294 214718 141326 214954
rect 141562 214718 141646 214954
rect 141882 214718 141914 214954
rect 141294 214634 141914 214718
rect 141294 214398 141326 214634
rect 141562 214398 141646 214634
rect 141882 214398 141914 214634
rect 141294 178954 141914 214398
rect 141294 178718 141326 178954
rect 141562 178718 141646 178954
rect 141882 178718 141914 178954
rect 141294 178634 141914 178718
rect 141294 178398 141326 178634
rect 141562 178398 141646 178634
rect 141882 178398 141914 178634
rect 141294 142954 141914 178398
rect 141294 142718 141326 142954
rect 141562 142718 141646 142954
rect 141882 142718 141914 142954
rect 141294 142634 141914 142718
rect 141294 142398 141326 142634
rect 141562 142398 141646 142634
rect 141882 142398 141914 142634
rect 141294 106954 141914 142398
rect 141294 106718 141326 106954
rect 141562 106718 141646 106954
rect 141882 106718 141914 106954
rect 141294 106634 141914 106718
rect 141294 106398 141326 106634
rect 141562 106398 141646 106634
rect 141882 106398 141914 106634
rect 141294 70954 141914 106398
rect 141294 70718 141326 70954
rect 141562 70718 141646 70954
rect 141882 70718 141914 70954
rect 141294 70634 141914 70718
rect 141294 70398 141326 70634
rect 141562 70398 141646 70634
rect 141882 70398 141914 70634
rect 141294 34954 141914 70398
rect 141294 34718 141326 34954
rect 141562 34718 141646 34954
rect 141882 34718 141914 34954
rect 141294 34634 141914 34718
rect 141294 34398 141326 34634
rect 141562 34398 141646 34634
rect 141882 34398 141914 34634
rect 141294 -7066 141914 34398
rect 141294 -7302 141326 -7066
rect 141562 -7302 141646 -7066
rect 141882 -7302 141914 -7066
rect 141294 -7386 141914 -7302
rect 141294 -7622 141326 -7386
rect 141562 -7622 141646 -7386
rect 141882 -7622 141914 -7386
rect 141294 -7654 141914 -7622
rect 145794 471454 146414 498000
rect 145794 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 146414 471454
rect 145794 471134 146414 471218
rect 145794 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 146414 471134
rect 145794 435454 146414 470898
rect 145794 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 146414 435454
rect 145794 435134 146414 435218
rect 145794 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 146414 435134
rect 145794 399454 146414 434898
rect 145794 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 146414 399454
rect 145794 399134 146414 399218
rect 145794 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 146414 399134
rect 145794 363454 146414 398898
rect 145794 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 146414 363454
rect 145794 363134 146414 363218
rect 145794 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 146414 363134
rect 145794 327454 146414 362898
rect 145794 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 146414 327454
rect 145794 327134 146414 327218
rect 145794 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 146414 327134
rect 145794 291454 146414 326898
rect 145794 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 146414 291454
rect 145794 291134 146414 291218
rect 145794 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 146414 291134
rect 145794 255454 146414 290898
rect 145794 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 146414 255454
rect 145794 255134 146414 255218
rect 145794 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 146414 255134
rect 145794 219454 146414 254898
rect 145794 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 146414 219454
rect 145794 219134 146414 219218
rect 145794 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 146414 219134
rect 145794 183454 146414 218898
rect 145794 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 146414 183454
rect 145794 183134 146414 183218
rect 145794 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 146414 183134
rect 145794 147454 146414 182898
rect 145794 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 146414 147454
rect 145794 147134 146414 147218
rect 145794 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 146414 147134
rect 145794 111454 146414 146898
rect 145794 111218 145826 111454
rect 146062 111218 146146 111454
rect 146382 111218 146414 111454
rect 145794 111134 146414 111218
rect 145794 110898 145826 111134
rect 146062 110898 146146 111134
rect 146382 110898 146414 111134
rect 145794 75454 146414 110898
rect 145794 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 146414 75454
rect 145794 75134 146414 75218
rect 145794 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 146414 75134
rect 145794 39454 146414 74898
rect 145794 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 146414 39454
rect 145794 39134 146414 39218
rect 145794 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 146414 39134
rect 145794 3454 146414 38898
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -7654 146414 -902
rect 150294 475954 150914 498000
rect 150294 475718 150326 475954
rect 150562 475718 150646 475954
rect 150882 475718 150914 475954
rect 150294 475634 150914 475718
rect 150294 475398 150326 475634
rect 150562 475398 150646 475634
rect 150882 475398 150914 475634
rect 150294 439954 150914 475398
rect 150294 439718 150326 439954
rect 150562 439718 150646 439954
rect 150882 439718 150914 439954
rect 150294 439634 150914 439718
rect 150294 439398 150326 439634
rect 150562 439398 150646 439634
rect 150882 439398 150914 439634
rect 150294 403954 150914 439398
rect 150294 403718 150326 403954
rect 150562 403718 150646 403954
rect 150882 403718 150914 403954
rect 150294 403634 150914 403718
rect 150294 403398 150326 403634
rect 150562 403398 150646 403634
rect 150882 403398 150914 403634
rect 150294 367954 150914 403398
rect 150294 367718 150326 367954
rect 150562 367718 150646 367954
rect 150882 367718 150914 367954
rect 150294 367634 150914 367718
rect 150294 367398 150326 367634
rect 150562 367398 150646 367634
rect 150882 367398 150914 367634
rect 150294 331954 150914 367398
rect 150294 331718 150326 331954
rect 150562 331718 150646 331954
rect 150882 331718 150914 331954
rect 150294 331634 150914 331718
rect 150294 331398 150326 331634
rect 150562 331398 150646 331634
rect 150882 331398 150914 331634
rect 150294 295954 150914 331398
rect 150294 295718 150326 295954
rect 150562 295718 150646 295954
rect 150882 295718 150914 295954
rect 150294 295634 150914 295718
rect 150294 295398 150326 295634
rect 150562 295398 150646 295634
rect 150882 295398 150914 295634
rect 150294 259954 150914 295398
rect 150294 259718 150326 259954
rect 150562 259718 150646 259954
rect 150882 259718 150914 259954
rect 150294 259634 150914 259718
rect 150294 259398 150326 259634
rect 150562 259398 150646 259634
rect 150882 259398 150914 259634
rect 150294 223954 150914 259398
rect 150294 223718 150326 223954
rect 150562 223718 150646 223954
rect 150882 223718 150914 223954
rect 150294 223634 150914 223718
rect 150294 223398 150326 223634
rect 150562 223398 150646 223634
rect 150882 223398 150914 223634
rect 150294 187954 150914 223398
rect 150294 187718 150326 187954
rect 150562 187718 150646 187954
rect 150882 187718 150914 187954
rect 150294 187634 150914 187718
rect 150294 187398 150326 187634
rect 150562 187398 150646 187634
rect 150882 187398 150914 187634
rect 150294 151954 150914 187398
rect 150294 151718 150326 151954
rect 150562 151718 150646 151954
rect 150882 151718 150914 151954
rect 150294 151634 150914 151718
rect 150294 151398 150326 151634
rect 150562 151398 150646 151634
rect 150882 151398 150914 151634
rect 150294 115954 150914 151398
rect 150294 115718 150326 115954
rect 150562 115718 150646 115954
rect 150882 115718 150914 115954
rect 150294 115634 150914 115718
rect 150294 115398 150326 115634
rect 150562 115398 150646 115634
rect 150882 115398 150914 115634
rect 150294 79954 150914 115398
rect 150294 79718 150326 79954
rect 150562 79718 150646 79954
rect 150882 79718 150914 79954
rect 150294 79634 150914 79718
rect 150294 79398 150326 79634
rect 150562 79398 150646 79634
rect 150882 79398 150914 79634
rect 150294 43954 150914 79398
rect 150294 43718 150326 43954
rect 150562 43718 150646 43954
rect 150882 43718 150914 43954
rect 150294 43634 150914 43718
rect 150294 43398 150326 43634
rect 150562 43398 150646 43634
rect 150882 43398 150914 43634
rect 150294 7954 150914 43398
rect 150294 7718 150326 7954
rect 150562 7718 150646 7954
rect 150882 7718 150914 7954
rect 150294 7634 150914 7718
rect 150294 7398 150326 7634
rect 150562 7398 150646 7634
rect 150882 7398 150914 7634
rect 150294 -1306 150914 7398
rect 150294 -1542 150326 -1306
rect 150562 -1542 150646 -1306
rect 150882 -1542 150914 -1306
rect 150294 -1626 150914 -1542
rect 150294 -1862 150326 -1626
rect 150562 -1862 150646 -1626
rect 150882 -1862 150914 -1626
rect 150294 -7654 150914 -1862
rect 154794 480454 155414 498000
rect 155542 496909 155602 499530
rect 160510 499530 160588 499590
rect 155539 496908 155605 496909
rect 155539 496844 155540 496908
rect 155604 496844 155605 496908
rect 155539 496843 155605 496844
rect 154794 480218 154826 480454
rect 155062 480218 155146 480454
rect 155382 480218 155414 480454
rect 154794 480134 155414 480218
rect 154794 479898 154826 480134
rect 155062 479898 155146 480134
rect 155382 479898 155414 480134
rect 154794 444454 155414 479898
rect 154794 444218 154826 444454
rect 155062 444218 155146 444454
rect 155382 444218 155414 444454
rect 154794 444134 155414 444218
rect 154794 443898 154826 444134
rect 155062 443898 155146 444134
rect 155382 443898 155414 444134
rect 154794 408454 155414 443898
rect 154794 408218 154826 408454
rect 155062 408218 155146 408454
rect 155382 408218 155414 408454
rect 154794 408134 155414 408218
rect 154794 407898 154826 408134
rect 155062 407898 155146 408134
rect 155382 407898 155414 408134
rect 154794 372454 155414 407898
rect 154794 372218 154826 372454
rect 155062 372218 155146 372454
rect 155382 372218 155414 372454
rect 154794 372134 155414 372218
rect 154794 371898 154826 372134
rect 155062 371898 155146 372134
rect 155382 371898 155414 372134
rect 154794 336454 155414 371898
rect 154794 336218 154826 336454
rect 155062 336218 155146 336454
rect 155382 336218 155414 336454
rect 154794 336134 155414 336218
rect 154794 335898 154826 336134
rect 155062 335898 155146 336134
rect 155382 335898 155414 336134
rect 154794 300454 155414 335898
rect 154794 300218 154826 300454
rect 155062 300218 155146 300454
rect 155382 300218 155414 300454
rect 154794 300134 155414 300218
rect 154794 299898 154826 300134
rect 155062 299898 155146 300134
rect 155382 299898 155414 300134
rect 154794 264454 155414 299898
rect 154794 264218 154826 264454
rect 155062 264218 155146 264454
rect 155382 264218 155414 264454
rect 154794 264134 155414 264218
rect 154794 263898 154826 264134
rect 155062 263898 155146 264134
rect 155382 263898 155414 264134
rect 154794 228454 155414 263898
rect 154794 228218 154826 228454
rect 155062 228218 155146 228454
rect 155382 228218 155414 228454
rect 154794 228134 155414 228218
rect 154794 227898 154826 228134
rect 155062 227898 155146 228134
rect 155382 227898 155414 228134
rect 154794 192454 155414 227898
rect 154794 192218 154826 192454
rect 155062 192218 155146 192454
rect 155382 192218 155414 192454
rect 154794 192134 155414 192218
rect 154794 191898 154826 192134
rect 155062 191898 155146 192134
rect 155382 191898 155414 192134
rect 154794 156454 155414 191898
rect 154794 156218 154826 156454
rect 155062 156218 155146 156454
rect 155382 156218 155414 156454
rect 154794 156134 155414 156218
rect 154794 155898 154826 156134
rect 155062 155898 155146 156134
rect 155382 155898 155414 156134
rect 154794 120454 155414 155898
rect 154794 120218 154826 120454
rect 155062 120218 155146 120454
rect 155382 120218 155414 120454
rect 154794 120134 155414 120218
rect 154794 119898 154826 120134
rect 155062 119898 155146 120134
rect 155382 119898 155414 120134
rect 154794 84454 155414 119898
rect 154794 84218 154826 84454
rect 155062 84218 155146 84454
rect 155382 84218 155414 84454
rect 154794 84134 155414 84218
rect 154794 83898 154826 84134
rect 155062 83898 155146 84134
rect 155382 83898 155414 84134
rect 154794 48454 155414 83898
rect 154794 48218 154826 48454
rect 155062 48218 155146 48454
rect 155382 48218 155414 48454
rect 154794 48134 155414 48218
rect 154794 47898 154826 48134
rect 155062 47898 155146 48134
rect 155382 47898 155414 48134
rect 154794 12454 155414 47898
rect 154794 12218 154826 12454
rect 155062 12218 155146 12454
rect 155382 12218 155414 12454
rect 154794 12134 155414 12218
rect 154794 11898 154826 12134
rect 155062 11898 155146 12134
rect 155382 11898 155414 12134
rect 154794 -2266 155414 11898
rect 154794 -2502 154826 -2266
rect 155062 -2502 155146 -2266
rect 155382 -2502 155414 -2266
rect 154794 -2586 155414 -2502
rect 154794 -2822 154826 -2586
rect 155062 -2822 155146 -2586
rect 155382 -2822 155414 -2586
rect 154794 -7654 155414 -2822
rect 159294 484954 159914 498000
rect 160510 496909 160570 499530
rect 160507 496908 160573 496909
rect 160507 496844 160508 496908
rect 160572 496844 160573 496908
rect 160507 496843 160573 496844
rect 159294 484718 159326 484954
rect 159562 484718 159646 484954
rect 159882 484718 159914 484954
rect 159294 484634 159914 484718
rect 159294 484398 159326 484634
rect 159562 484398 159646 484634
rect 159882 484398 159914 484634
rect 159294 448954 159914 484398
rect 159294 448718 159326 448954
rect 159562 448718 159646 448954
rect 159882 448718 159914 448954
rect 159294 448634 159914 448718
rect 159294 448398 159326 448634
rect 159562 448398 159646 448634
rect 159882 448398 159914 448634
rect 159294 412954 159914 448398
rect 159294 412718 159326 412954
rect 159562 412718 159646 412954
rect 159882 412718 159914 412954
rect 159294 412634 159914 412718
rect 159294 412398 159326 412634
rect 159562 412398 159646 412634
rect 159882 412398 159914 412634
rect 159294 376954 159914 412398
rect 159294 376718 159326 376954
rect 159562 376718 159646 376954
rect 159882 376718 159914 376954
rect 159294 376634 159914 376718
rect 159294 376398 159326 376634
rect 159562 376398 159646 376634
rect 159882 376398 159914 376634
rect 159294 340954 159914 376398
rect 159294 340718 159326 340954
rect 159562 340718 159646 340954
rect 159882 340718 159914 340954
rect 159294 340634 159914 340718
rect 159294 340398 159326 340634
rect 159562 340398 159646 340634
rect 159882 340398 159914 340634
rect 159294 304954 159914 340398
rect 159294 304718 159326 304954
rect 159562 304718 159646 304954
rect 159882 304718 159914 304954
rect 159294 304634 159914 304718
rect 159294 304398 159326 304634
rect 159562 304398 159646 304634
rect 159882 304398 159914 304634
rect 159294 268954 159914 304398
rect 159294 268718 159326 268954
rect 159562 268718 159646 268954
rect 159882 268718 159914 268954
rect 159294 268634 159914 268718
rect 159294 268398 159326 268634
rect 159562 268398 159646 268634
rect 159882 268398 159914 268634
rect 159294 232954 159914 268398
rect 159294 232718 159326 232954
rect 159562 232718 159646 232954
rect 159882 232718 159914 232954
rect 159294 232634 159914 232718
rect 159294 232398 159326 232634
rect 159562 232398 159646 232634
rect 159882 232398 159914 232634
rect 159294 196954 159914 232398
rect 159294 196718 159326 196954
rect 159562 196718 159646 196954
rect 159882 196718 159914 196954
rect 159294 196634 159914 196718
rect 159294 196398 159326 196634
rect 159562 196398 159646 196634
rect 159882 196398 159914 196634
rect 159294 160954 159914 196398
rect 159294 160718 159326 160954
rect 159562 160718 159646 160954
rect 159882 160718 159914 160954
rect 159294 160634 159914 160718
rect 159294 160398 159326 160634
rect 159562 160398 159646 160634
rect 159882 160398 159914 160634
rect 159294 124954 159914 160398
rect 159294 124718 159326 124954
rect 159562 124718 159646 124954
rect 159882 124718 159914 124954
rect 159294 124634 159914 124718
rect 159294 124398 159326 124634
rect 159562 124398 159646 124634
rect 159882 124398 159914 124634
rect 159294 88954 159914 124398
rect 159294 88718 159326 88954
rect 159562 88718 159646 88954
rect 159882 88718 159914 88954
rect 159294 88634 159914 88718
rect 159294 88398 159326 88634
rect 159562 88398 159646 88634
rect 159882 88398 159914 88634
rect 159294 52954 159914 88398
rect 159294 52718 159326 52954
rect 159562 52718 159646 52954
rect 159882 52718 159914 52954
rect 159294 52634 159914 52718
rect 159294 52398 159326 52634
rect 159562 52398 159646 52634
rect 159882 52398 159914 52634
rect 159294 16954 159914 52398
rect 159294 16718 159326 16954
rect 159562 16718 159646 16954
rect 159882 16718 159914 16954
rect 159294 16634 159914 16718
rect 159294 16398 159326 16634
rect 159562 16398 159646 16634
rect 159882 16398 159914 16634
rect 159294 -3226 159914 16398
rect 159294 -3462 159326 -3226
rect 159562 -3462 159646 -3226
rect 159882 -3462 159914 -3226
rect 159294 -3546 159914 -3462
rect 159294 -3782 159326 -3546
rect 159562 -3782 159646 -3546
rect 159882 -3782 159914 -3546
rect 159294 -7654 159914 -3782
rect 163794 489454 164414 498000
rect 163794 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 164414 489454
rect 163794 489134 164414 489218
rect 163794 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 164414 489134
rect 163794 453454 164414 488898
rect 163794 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 164414 453454
rect 163794 453134 164414 453218
rect 163794 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 164414 453134
rect 163794 417454 164414 452898
rect 163794 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 164414 417454
rect 163794 417134 164414 417218
rect 163794 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 164414 417134
rect 163794 381454 164414 416898
rect 163794 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 164414 381454
rect 163794 381134 164414 381218
rect 163794 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 164414 381134
rect 163794 345454 164414 380898
rect 163794 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 164414 345454
rect 163794 345134 164414 345218
rect 163794 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 164414 345134
rect 163794 309454 164414 344898
rect 163794 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 164414 309454
rect 163794 309134 164414 309218
rect 163794 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 164414 309134
rect 163794 273454 164414 308898
rect 163794 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 164414 273454
rect 163794 273134 164414 273218
rect 163794 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 164414 273134
rect 163794 237454 164414 272898
rect 163794 237218 163826 237454
rect 164062 237218 164146 237454
rect 164382 237218 164414 237454
rect 163794 237134 164414 237218
rect 163794 236898 163826 237134
rect 164062 236898 164146 237134
rect 164382 236898 164414 237134
rect 163794 201454 164414 236898
rect 163794 201218 163826 201454
rect 164062 201218 164146 201454
rect 164382 201218 164414 201454
rect 163794 201134 164414 201218
rect 163794 200898 163826 201134
rect 164062 200898 164146 201134
rect 164382 200898 164414 201134
rect 163794 165454 164414 200898
rect 163794 165218 163826 165454
rect 164062 165218 164146 165454
rect 164382 165218 164414 165454
rect 163794 165134 164414 165218
rect 163794 164898 163826 165134
rect 164062 164898 164146 165134
rect 164382 164898 164414 165134
rect 163794 129454 164414 164898
rect 163794 129218 163826 129454
rect 164062 129218 164146 129454
rect 164382 129218 164414 129454
rect 163794 129134 164414 129218
rect 163794 128898 163826 129134
rect 164062 128898 164146 129134
rect 164382 128898 164414 129134
rect 163794 93454 164414 128898
rect 163794 93218 163826 93454
rect 164062 93218 164146 93454
rect 164382 93218 164414 93454
rect 163794 93134 164414 93218
rect 163794 92898 163826 93134
rect 164062 92898 164146 93134
rect 164382 92898 164414 93134
rect 163794 57454 164414 92898
rect 163794 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 164414 57454
rect 163794 57134 164414 57218
rect 163794 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 164414 57134
rect 163794 21454 164414 56898
rect 163794 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 164414 21454
rect 163794 21134 164414 21218
rect 163794 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 164414 21134
rect 163794 -4186 164414 20898
rect 163794 -4422 163826 -4186
rect 164062 -4422 164146 -4186
rect 164382 -4422 164414 -4186
rect 163794 -4506 164414 -4422
rect 163794 -4742 163826 -4506
rect 164062 -4742 164146 -4506
rect 164382 -4742 164414 -4506
rect 163794 -7654 164414 -4742
rect 168294 493954 168914 498000
rect 168294 493718 168326 493954
rect 168562 493718 168646 493954
rect 168882 493718 168914 493954
rect 168294 493634 168914 493718
rect 168294 493398 168326 493634
rect 168562 493398 168646 493634
rect 168882 493398 168914 493634
rect 168294 457954 168914 493398
rect 168294 457718 168326 457954
rect 168562 457718 168646 457954
rect 168882 457718 168914 457954
rect 168294 457634 168914 457718
rect 168294 457398 168326 457634
rect 168562 457398 168646 457634
rect 168882 457398 168914 457634
rect 168294 421954 168914 457398
rect 168294 421718 168326 421954
rect 168562 421718 168646 421954
rect 168882 421718 168914 421954
rect 168294 421634 168914 421718
rect 168294 421398 168326 421634
rect 168562 421398 168646 421634
rect 168882 421398 168914 421634
rect 168294 385954 168914 421398
rect 168294 385718 168326 385954
rect 168562 385718 168646 385954
rect 168882 385718 168914 385954
rect 168294 385634 168914 385718
rect 168294 385398 168326 385634
rect 168562 385398 168646 385634
rect 168882 385398 168914 385634
rect 168294 349954 168914 385398
rect 168294 349718 168326 349954
rect 168562 349718 168646 349954
rect 168882 349718 168914 349954
rect 168294 349634 168914 349718
rect 168294 349398 168326 349634
rect 168562 349398 168646 349634
rect 168882 349398 168914 349634
rect 168294 313954 168914 349398
rect 168294 313718 168326 313954
rect 168562 313718 168646 313954
rect 168882 313718 168914 313954
rect 168294 313634 168914 313718
rect 168294 313398 168326 313634
rect 168562 313398 168646 313634
rect 168882 313398 168914 313634
rect 168294 277954 168914 313398
rect 168294 277718 168326 277954
rect 168562 277718 168646 277954
rect 168882 277718 168914 277954
rect 168294 277634 168914 277718
rect 168294 277398 168326 277634
rect 168562 277398 168646 277634
rect 168882 277398 168914 277634
rect 168294 241954 168914 277398
rect 168294 241718 168326 241954
rect 168562 241718 168646 241954
rect 168882 241718 168914 241954
rect 168294 241634 168914 241718
rect 168294 241398 168326 241634
rect 168562 241398 168646 241634
rect 168882 241398 168914 241634
rect 168294 205954 168914 241398
rect 168294 205718 168326 205954
rect 168562 205718 168646 205954
rect 168882 205718 168914 205954
rect 168294 205634 168914 205718
rect 168294 205398 168326 205634
rect 168562 205398 168646 205634
rect 168882 205398 168914 205634
rect 168294 169954 168914 205398
rect 168294 169718 168326 169954
rect 168562 169718 168646 169954
rect 168882 169718 168914 169954
rect 168294 169634 168914 169718
rect 168294 169398 168326 169634
rect 168562 169398 168646 169634
rect 168882 169398 168914 169634
rect 168294 133954 168914 169398
rect 168294 133718 168326 133954
rect 168562 133718 168646 133954
rect 168882 133718 168914 133954
rect 168294 133634 168914 133718
rect 168294 133398 168326 133634
rect 168562 133398 168646 133634
rect 168882 133398 168914 133634
rect 168294 97954 168914 133398
rect 168294 97718 168326 97954
rect 168562 97718 168646 97954
rect 168882 97718 168914 97954
rect 168294 97634 168914 97718
rect 168294 97398 168326 97634
rect 168562 97398 168646 97634
rect 168882 97398 168914 97634
rect 168294 61954 168914 97398
rect 168294 61718 168326 61954
rect 168562 61718 168646 61954
rect 168882 61718 168914 61954
rect 168294 61634 168914 61718
rect 168294 61398 168326 61634
rect 168562 61398 168646 61634
rect 168882 61398 168914 61634
rect 168294 25954 168914 61398
rect 168294 25718 168326 25954
rect 168562 25718 168646 25954
rect 168882 25718 168914 25954
rect 168294 25634 168914 25718
rect 168294 25398 168326 25634
rect 168562 25398 168646 25634
rect 168882 25398 168914 25634
rect 168294 -5146 168914 25398
rect 168294 -5382 168326 -5146
rect 168562 -5382 168646 -5146
rect 168882 -5382 168914 -5146
rect 168294 -5466 168914 -5382
rect 168294 -5702 168326 -5466
rect 168562 -5702 168646 -5466
rect 168882 -5702 168914 -5466
rect 168294 -7654 168914 -5702
rect 172794 462454 173414 498000
rect 172794 462218 172826 462454
rect 173062 462218 173146 462454
rect 173382 462218 173414 462454
rect 172794 462134 173414 462218
rect 172794 461898 172826 462134
rect 173062 461898 173146 462134
rect 173382 461898 173414 462134
rect 172794 426454 173414 461898
rect 172794 426218 172826 426454
rect 173062 426218 173146 426454
rect 173382 426218 173414 426454
rect 172794 426134 173414 426218
rect 172794 425898 172826 426134
rect 173062 425898 173146 426134
rect 173382 425898 173414 426134
rect 172794 390454 173414 425898
rect 172794 390218 172826 390454
rect 173062 390218 173146 390454
rect 173382 390218 173414 390454
rect 172794 390134 173414 390218
rect 172794 389898 172826 390134
rect 173062 389898 173146 390134
rect 173382 389898 173414 390134
rect 172794 354454 173414 389898
rect 172794 354218 172826 354454
rect 173062 354218 173146 354454
rect 173382 354218 173414 354454
rect 172794 354134 173414 354218
rect 172794 353898 172826 354134
rect 173062 353898 173146 354134
rect 173382 353898 173414 354134
rect 172794 318454 173414 353898
rect 172794 318218 172826 318454
rect 173062 318218 173146 318454
rect 173382 318218 173414 318454
rect 172794 318134 173414 318218
rect 172794 317898 172826 318134
rect 173062 317898 173146 318134
rect 173382 317898 173414 318134
rect 172794 282454 173414 317898
rect 172794 282218 172826 282454
rect 173062 282218 173146 282454
rect 173382 282218 173414 282454
rect 172794 282134 173414 282218
rect 172794 281898 172826 282134
rect 173062 281898 173146 282134
rect 173382 281898 173414 282134
rect 172794 246454 173414 281898
rect 172794 246218 172826 246454
rect 173062 246218 173146 246454
rect 173382 246218 173414 246454
rect 172794 246134 173414 246218
rect 172794 245898 172826 246134
rect 173062 245898 173146 246134
rect 173382 245898 173414 246134
rect 172794 210454 173414 245898
rect 172794 210218 172826 210454
rect 173062 210218 173146 210454
rect 173382 210218 173414 210454
rect 172794 210134 173414 210218
rect 172794 209898 172826 210134
rect 173062 209898 173146 210134
rect 173382 209898 173414 210134
rect 172794 174454 173414 209898
rect 172794 174218 172826 174454
rect 173062 174218 173146 174454
rect 173382 174218 173414 174454
rect 172794 174134 173414 174218
rect 172794 173898 172826 174134
rect 173062 173898 173146 174134
rect 173382 173898 173414 174134
rect 172794 138454 173414 173898
rect 172794 138218 172826 138454
rect 173062 138218 173146 138454
rect 173382 138218 173414 138454
rect 172794 138134 173414 138218
rect 172794 137898 172826 138134
rect 173062 137898 173146 138134
rect 173382 137898 173414 138134
rect 172794 102454 173414 137898
rect 172794 102218 172826 102454
rect 173062 102218 173146 102454
rect 173382 102218 173414 102454
rect 172794 102134 173414 102218
rect 172794 101898 172826 102134
rect 173062 101898 173146 102134
rect 173382 101898 173414 102134
rect 172794 66454 173414 101898
rect 172794 66218 172826 66454
rect 173062 66218 173146 66454
rect 173382 66218 173414 66454
rect 172794 66134 173414 66218
rect 172794 65898 172826 66134
rect 173062 65898 173146 66134
rect 173382 65898 173414 66134
rect 172794 30454 173414 65898
rect 172794 30218 172826 30454
rect 173062 30218 173146 30454
rect 173382 30218 173414 30454
rect 172794 30134 173414 30218
rect 172794 29898 172826 30134
rect 173062 29898 173146 30134
rect 173382 29898 173414 30134
rect 172794 -6106 173414 29898
rect 172794 -6342 172826 -6106
rect 173062 -6342 173146 -6106
rect 173382 -6342 173414 -6106
rect 172794 -6426 173414 -6342
rect 172794 -6662 172826 -6426
rect 173062 -6662 173146 -6426
rect 173382 -6662 173414 -6426
rect 172794 -7654 173414 -6662
rect 177294 466954 177914 498000
rect 177294 466718 177326 466954
rect 177562 466718 177646 466954
rect 177882 466718 177914 466954
rect 177294 466634 177914 466718
rect 177294 466398 177326 466634
rect 177562 466398 177646 466634
rect 177882 466398 177914 466634
rect 177294 430954 177914 466398
rect 177294 430718 177326 430954
rect 177562 430718 177646 430954
rect 177882 430718 177914 430954
rect 177294 430634 177914 430718
rect 177294 430398 177326 430634
rect 177562 430398 177646 430634
rect 177882 430398 177914 430634
rect 177294 394954 177914 430398
rect 177294 394718 177326 394954
rect 177562 394718 177646 394954
rect 177882 394718 177914 394954
rect 177294 394634 177914 394718
rect 177294 394398 177326 394634
rect 177562 394398 177646 394634
rect 177882 394398 177914 394634
rect 177294 358954 177914 394398
rect 177294 358718 177326 358954
rect 177562 358718 177646 358954
rect 177882 358718 177914 358954
rect 177294 358634 177914 358718
rect 177294 358398 177326 358634
rect 177562 358398 177646 358634
rect 177882 358398 177914 358634
rect 177294 322954 177914 358398
rect 177294 322718 177326 322954
rect 177562 322718 177646 322954
rect 177882 322718 177914 322954
rect 177294 322634 177914 322718
rect 177294 322398 177326 322634
rect 177562 322398 177646 322634
rect 177882 322398 177914 322634
rect 177294 286954 177914 322398
rect 177294 286718 177326 286954
rect 177562 286718 177646 286954
rect 177882 286718 177914 286954
rect 177294 286634 177914 286718
rect 177294 286398 177326 286634
rect 177562 286398 177646 286634
rect 177882 286398 177914 286634
rect 177294 250954 177914 286398
rect 177294 250718 177326 250954
rect 177562 250718 177646 250954
rect 177882 250718 177914 250954
rect 177294 250634 177914 250718
rect 177294 250398 177326 250634
rect 177562 250398 177646 250634
rect 177882 250398 177914 250634
rect 177294 214954 177914 250398
rect 177294 214718 177326 214954
rect 177562 214718 177646 214954
rect 177882 214718 177914 214954
rect 177294 214634 177914 214718
rect 177294 214398 177326 214634
rect 177562 214398 177646 214634
rect 177882 214398 177914 214634
rect 177294 178954 177914 214398
rect 177294 178718 177326 178954
rect 177562 178718 177646 178954
rect 177882 178718 177914 178954
rect 177294 178634 177914 178718
rect 177294 178398 177326 178634
rect 177562 178398 177646 178634
rect 177882 178398 177914 178634
rect 177294 142954 177914 178398
rect 177294 142718 177326 142954
rect 177562 142718 177646 142954
rect 177882 142718 177914 142954
rect 177294 142634 177914 142718
rect 177294 142398 177326 142634
rect 177562 142398 177646 142634
rect 177882 142398 177914 142634
rect 177294 106954 177914 142398
rect 177294 106718 177326 106954
rect 177562 106718 177646 106954
rect 177882 106718 177914 106954
rect 177294 106634 177914 106718
rect 177294 106398 177326 106634
rect 177562 106398 177646 106634
rect 177882 106398 177914 106634
rect 177294 70954 177914 106398
rect 177294 70718 177326 70954
rect 177562 70718 177646 70954
rect 177882 70718 177914 70954
rect 177294 70634 177914 70718
rect 177294 70398 177326 70634
rect 177562 70398 177646 70634
rect 177882 70398 177914 70634
rect 177294 34954 177914 70398
rect 177294 34718 177326 34954
rect 177562 34718 177646 34954
rect 177882 34718 177914 34954
rect 177294 34634 177914 34718
rect 177294 34398 177326 34634
rect 177562 34398 177646 34634
rect 177882 34398 177914 34634
rect 177294 -7066 177914 34398
rect 177294 -7302 177326 -7066
rect 177562 -7302 177646 -7066
rect 177882 -7302 177914 -7066
rect 177294 -7386 177914 -7302
rect 177294 -7622 177326 -7386
rect 177562 -7622 177646 -7386
rect 177882 -7622 177914 -7386
rect 177294 -7654 177914 -7622
rect 181794 471454 182414 498000
rect 181794 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 182414 471454
rect 181794 471134 182414 471218
rect 181794 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 182414 471134
rect 181794 435454 182414 470898
rect 181794 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 182414 435454
rect 181794 435134 182414 435218
rect 181794 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 182414 435134
rect 181794 399454 182414 434898
rect 181794 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 182414 399454
rect 181794 399134 182414 399218
rect 181794 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 182414 399134
rect 181794 363454 182414 398898
rect 181794 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 182414 363454
rect 181794 363134 182414 363218
rect 181794 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 182414 363134
rect 181794 327454 182414 362898
rect 181794 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 182414 327454
rect 181794 327134 182414 327218
rect 181794 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 182414 327134
rect 181794 291454 182414 326898
rect 181794 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 182414 291454
rect 181794 291134 182414 291218
rect 181794 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 182414 291134
rect 181794 255454 182414 290898
rect 181794 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 182414 255454
rect 181794 255134 182414 255218
rect 181794 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 182414 255134
rect 181794 219454 182414 254898
rect 181794 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 182414 219454
rect 181794 219134 182414 219218
rect 181794 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 182414 219134
rect 181794 183454 182414 218898
rect 181794 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 182414 183454
rect 181794 183134 182414 183218
rect 181794 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 182414 183134
rect 181794 147454 182414 182898
rect 181794 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 182414 147454
rect 181794 147134 182414 147218
rect 181794 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 182414 147134
rect 181794 111454 182414 146898
rect 181794 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 182414 111454
rect 181794 111134 182414 111218
rect 181794 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 182414 111134
rect 181794 75454 182414 110898
rect 181794 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 182414 75454
rect 181794 75134 182414 75218
rect 181794 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 182414 75134
rect 181794 39454 182414 74898
rect 181794 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 182414 39454
rect 181794 39134 182414 39218
rect 181794 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 182414 39134
rect 181794 3454 182414 38898
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -7654 182414 -902
rect 186294 475954 186914 498000
rect 186294 475718 186326 475954
rect 186562 475718 186646 475954
rect 186882 475718 186914 475954
rect 186294 475634 186914 475718
rect 186294 475398 186326 475634
rect 186562 475398 186646 475634
rect 186882 475398 186914 475634
rect 186294 439954 186914 475398
rect 186294 439718 186326 439954
rect 186562 439718 186646 439954
rect 186882 439718 186914 439954
rect 186294 439634 186914 439718
rect 186294 439398 186326 439634
rect 186562 439398 186646 439634
rect 186882 439398 186914 439634
rect 186294 403954 186914 439398
rect 186294 403718 186326 403954
rect 186562 403718 186646 403954
rect 186882 403718 186914 403954
rect 186294 403634 186914 403718
rect 186294 403398 186326 403634
rect 186562 403398 186646 403634
rect 186882 403398 186914 403634
rect 186294 367954 186914 403398
rect 186294 367718 186326 367954
rect 186562 367718 186646 367954
rect 186882 367718 186914 367954
rect 186294 367634 186914 367718
rect 186294 367398 186326 367634
rect 186562 367398 186646 367634
rect 186882 367398 186914 367634
rect 186294 331954 186914 367398
rect 186294 331718 186326 331954
rect 186562 331718 186646 331954
rect 186882 331718 186914 331954
rect 186294 331634 186914 331718
rect 186294 331398 186326 331634
rect 186562 331398 186646 331634
rect 186882 331398 186914 331634
rect 186294 295954 186914 331398
rect 186294 295718 186326 295954
rect 186562 295718 186646 295954
rect 186882 295718 186914 295954
rect 186294 295634 186914 295718
rect 186294 295398 186326 295634
rect 186562 295398 186646 295634
rect 186882 295398 186914 295634
rect 186294 259954 186914 295398
rect 186294 259718 186326 259954
rect 186562 259718 186646 259954
rect 186882 259718 186914 259954
rect 186294 259634 186914 259718
rect 186294 259398 186326 259634
rect 186562 259398 186646 259634
rect 186882 259398 186914 259634
rect 186294 223954 186914 259398
rect 186294 223718 186326 223954
rect 186562 223718 186646 223954
rect 186882 223718 186914 223954
rect 186294 223634 186914 223718
rect 186294 223398 186326 223634
rect 186562 223398 186646 223634
rect 186882 223398 186914 223634
rect 186294 187954 186914 223398
rect 186294 187718 186326 187954
rect 186562 187718 186646 187954
rect 186882 187718 186914 187954
rect 186294 187634 186914 187718
rect 186294 187398 186326 187634
rect 186562 187398 186646 187634
rect 186882 187398 186914 187634
rect 186294 151954 186914 187398
rect 186294 151718 186326 151954
rect 186562 151718 186646 151954
rect 186882 151718 186914 151954
rect 186294 151634 186914 151718
rect 186294 151398 186326 151634
rect 186562 151398 186646 151634
rect 186882 151398 186914 151634
rect 186294 115954 186914 151398
rect 186294 115718 186326 115954
rect 186562 115718 186646 115954
rect 186882 115718 186914 115954
rect 186294 115634 186914 115718
rect 186294 115398 186326 115634
rect 186562 115398 186646 115634
rect 186882 115398 186914 115634
rect 186294 79954 186914 115398
rect 186294 79718 186326 79954
rect 186562 79718 186646 79954
rect 186882 79718 186914 79954
rect 186294 79634 186914 79718
rect 186294 79398 186326 79634
rect 186562 79398 186646 79634
rect 186882 79398 186914 79634
rect 186294 43954 186914 79398
rect 186294 43718 186326 43954
rect 186562 43718 186646 43954
rect 186882 43718 186914 43954
rect 186294 43634 186914 43718
rect 186294 43398 186326 43634
rect 186562 43398 186646 43634
rect 186882 43398 186914 43634
rect 186294 7954 186914 43398
rect 186294 7718 186326 7954
rect 186562 7718 186646 7954
rect 186882 7718 186914 7954
rect 186294 7634 186914 7718
rect 186294 7398 186326 7634
rect 186562 7398 186646 7634
rect 186882 7398 186914 7634
rect 186294 -1306 186914 7398
rect 186294 -1542 186326 -1306
rect 186562 -1542 186646 -1306
rect 186882 -1542 186914 -1306
rect 186294 -1626 186914 -1542
rect 186294 -1862 186326 -1626
rect 186562 -1862 186646 -1626
rect 186882 -1862 186914 -1626
rect 186294 -7654 186914 -1862
rect 190794 480454 191414 498000
rect 190794 480218 190826 480454
rect 191062 480218 191146 480454
rect 191382 480218 191414 480454
rect 190794 480134 191414 480218
rect 190794 479898 190826 480134
rect 191062 479898 191146 480134
rect 191382 479898 191414 480134
rect 190794 444454 191414 479898
rect 190794 444218 190826 444454
rect 191062 444218 191146 444454
rect 191382 444218 191414 444454
rect 190794 444134 191414 444218
rect 190794 443898 190826 444134
rect 191062 443898 191146 444134
rect 191382 443898 191414 444134
rect 190794 408454 191414 443898
rect 190794 408218 190826 408454
rect 191062 408218 191146 408454
rect 191382 408218 191414 408454
rect 190794 408134 191414 408218
rect 190794 407898 190826 408134
rect 191062 407898 191146 408134
rect 191382 407898 191414 408134
rect 190794 372454 191414 407898
rect 190794 372218 190826 372454
rect 191062 372218 191146 372454
rect 191382 372218 191414 372454
rect 190794 372134 191414 372218
rect 190794 371898 190826 372134
rect 191062 371898 191146 372134
rect 191382 371898 191414 372134
rect 190794 336454 191414 371898
rect 190794 336218 190826 336454
rect 191062 336218 191146 336454
rect 191382 336218 191414 336454
rect 190794 336134 191414 336218
rect 190794 335898 190826 336134
rect 191062 335898 191146 336134
rect 191382 335898 191414 336134
rect 190794 300454 191414 335898
rect 190794 300218 190826 300454
rect 191062 300218 191146 300454
rect 191382 300218 191414 300454
rect 190794 300134 191414 300218
rect 190794 299898 190826 300134
rect 191062 299898 191146 300134
rect 191382 299898 191414 300134
rect 190794 264454 191414 299898
rect 190794 264218 190826 264454
rect 191062 264218 191146 264454
rect 191382 264218 191414 264454
rect 190794 264134 191414 264218
rect 190794 263898 190826 264134
rect 191062 263898 191146 264134
rect 191382 263898 191414 264134
rect 190794 228454 191414 263898
rect 190794 228218 190826 228454
rect 191062 228218 191146 228454
rect 191382 228218 191414 228454
rect 190794 228134 191414 228218
rect 190794 227898 190826 228134
rect 191062 227898 191146 228134
rect 191382 227898 191414 228134
rect 190794 192454 191414 227898
rect 190794 192218 190826 192454
rect 191062 192218 191146 192454
rect 191382 192218 191414 192454
rect 190794 192134 191414 192218
rect 190794 191898 190826 192134
rect 191062 191898 191146 192134
rect 191382 191898 191414 192134
rect 190794 156454 191414 191898
rect 190794 156218 190826 156454
rect 191062 156218 191146 156454
rect 191382 156218 191414 156454
rect 190794 156134 191414 156218
rect 190794 155898 190826 156134
rect 191062 155898 191146 156134
rect 191382 155898 191414 156134
rect 190794 120454 191414 155898
rect 190794 120218 190826 120454
rect 191062 120218 191146 120454
rect 191382 120218 191414 120454
rect 190794 120134 191414 120218
rect 190794 119898 190826 120134
rect 191062 119898 191146 120134
rect 191382 119898 191414 120134
rect 190794 84454 191414 119898
rect 190794 84218 190826 84454
rect 191062 84218 191146 84454
rect 191382 84218 191414 84454
rect 190794 84134 191414 84218
rect 190794 83898 190826 84134
rect 191062 83898 191146 84134
rect 191382 83898 191414 84134
rect 190794 48454 191414 83898
rect 190794 48218 190826 48454
rect 191062 48218 191146 48454
rect 191382 48218 191414 48454
rect 190794 48134 191414 48218
rect 190794 47898 190826 48134
rect 191062 47898 191146 48134
rect 191382 47898 191414 48134
rect 190794 12454 191414 47898
rect 190794 12218 190826 12454
rect 191062 12218 191146 12454
rect 191382 12218 191414 12454
rect 190794 12134 191414 12218
rect 190794 11898 190826 12134
rect 191062 11898 191146 12134
rect 191382 11898 191414 12134
rect 190794 -2266 191414 11898
rect 190794 -2502 190826 -2266
rect 191062 -2502 191146 -2266
rect 191382 -2502 191414 -2266
rect 190794 -2586 191414 -2502
rect 190794 -2822 190826 -2586
rect 191062 -2822 191146 -2586
rect 191382 -2822 191414 -2586
rect 190794 -7654 191414 -2822
rect 195294 484954 195914 520398
rect 195294 484718 195326 484954
rect 195562 484718 195646 484954
rect 195882 484718 195914 484954
rect 195294 484634 195914 484718
rect 195294 484398 195326 484634
rect 195562 484398 195646 484634
rect 195882 484398 195914 484634
rect 195294 448954 195914 484398
rect 195294 448718 195326 448954
rect 195562 448718 195646 448954
rect 195882 448718 195914 448954
rect 195294 448634 195914 448718
rect 195294 448398 195326 448634
rect 195562 448398 195646 448634
rect 195882 448398 195914 448634
rect 195294 412954 195914 448398
rect 195294 412718 195326 412954
rect 195562 412718 195646 412954
rect 195882 412718 195914 412954
rect 195294 412634 195914 412718
rect 195294 412398 195326 412634
rect 195562 412398 195646 412634
rect 195882 412398 195914 412634
rect 195294 376954 195914 412398
rect 195294 376718 195326 376954
rect 195562 376718 195646 376954
rect 195882 376718 195914 376954
rect 195294 376634 195914 376718
rect 195294 376398 195326 376634
rect 195562 376398 195646 376634
rect 195882 376398 195914 376634
rect 195294 340954 195914 376398
rect 195294 340718 195326 340954
rect 195562 340718 195646 340954
rect 195882 340718 195914 340954
rect 195294 340634 195914 340718
rect 195294 340398 195326 340634
rect 195562 340398 195646 340634
rect 195882 340398 195914 340634
rect 195294 304954 195914 340398
rect 195294 304718 195326 304954
rect 195562 304718 195646 304954
rect 195882 304718 195914 304954
rect 195294 304634 195914 304718
rect 195294 304398 195326 304634
rect 195562 304398 195646 304634
rect 195882 304398 195914 304634
rect 195294 268954 195914 304398
rect 195294 268718 195326 268954
rect 195562 268718 195646 268954
rect 195882 268718 195914 268954
rect 195294 268634 195914 268718
rect 195294 268398 195326 268634
rect 195562 268398 195646 268634
rect 195882 268398 195914 268634
rect 195294 232954 195914 268398
rect 195294 232718 195326 232954
rect 195562 232718 195646 232954
rect 195882 232718 195914 232954
rect 195294 232634 195914 232718
rect 195294 232398 195326 232634
rect 195562 232398 195646 232634
rect 195882 232398 195914 232634
rect 195294 196954 195914 232398
rect 195294 196718 195326 196954
rect 195562 196718 195646 196954
rect 195882 196718 195914 196954
rect 195294 196634 195914 196718
rect 195294 196398 195326 196634
rect 195562 196398 195646 196634
rect 195882 196398 195914 196634
rect 195294 160954 195914 196398
rect 195294 160718 195326 160954
rect 195562 160718 195646 160954
rect 195882 160718 195914 160954
rect 195294 160634 195914 160718
rect 195294 160398 195326 160634
rect 195562 160398 195646 160634
rect 195882 160398 195914 160634
rect 195294 124954 195914 160398
rect 195294 124718 195326 124954
rect 195562 124718 195646 124954
rect 195882 124718 195914 124954
rect 195294 124634 195914 124718
rect 195294 124398 195326 124634
rect 195562 124398 195646 124634
rect 195882 124398 195914 124634
rect 195294 88954 195914 124398
rect 195294 88718 195326 88954
rect 195562 88718 195646 88954
rect 195882 88718 195914 88954
rect 195294 88634 195914 88718
rect 195294 88398 195326 88634
rect 195562 88398 195646 88634
rect 195882 88398 195914 88634
rect 195294 52954 195914 88398
rect 195294 52718 195326 52954
rect 195562 52718 195646 52954
rect 195882 52718 195914 52954
rect 195294 52634 195914 52718
rect 195294 52398 195326 52634
rect 195562 52398 195646 52634
rect 195882 52398 195914 52634
rect 195294 16954 195914 52398
rect 195294 16718 195326 16954
rect 195562 16718 195646 16954
rect 195882 16718 195914 16954
rect 195294 16634 195914 16718
rect 195294 16398 195326 16634
rect 195562 16398 195646 16634
rect 195882 16398 195914 16634
rect 195294 -3226 195914 16398
rect 195294 -3462 195326 -3226
rect 195562 -3462 195646 -3226
rect 195882 -3462 195914 -3226
rect 195294 -3546 195914 -3462
rect 195294 -3782 195326 -3546
rect 195562 -3782 195646 -3546
rect 195882 -3782 195914 -3546
rect 195294 -7654 195914 -3782
rect 199794 708678 200414 711590
rect 199794 708442 199826 708678
rect 200062 708442 200146 708678
rect 200382 708442 200414 708678
rect 199794 708358 200414 708442
rect 199794 708122 199826 708358
rect 200062 708122 200146 708358
rect 200382 708122 200414 708358
rect 199794 669454 200414 708122
rect 199794 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 200414 669454
rect 199794 669134 200414 669218
rect 199794 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 200414 669134
rect 199794 633454 200414 668898
rect 199794 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 200414 633454
rect 199794 633134 200414 633218
rect 199794 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 200414 633134
rect 199794 597454 200414 632898
rect 199794 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 200414 597454
rect 199794 597134 200414 597218
rect 199794 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 200414 597134
rect 199794 561454 200414 596898
rect 199794 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 200414 561454
rect 199794 561134 200414 561218
rect 199794 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 200414 561134
rect 199794 525454 200414 560898
rect 199794 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 200414 525454
rect 199794 525134 200414 525218
rect 199794 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 200414 525134
rect 199794 489454 200414 524898
rect 199794 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 200414 489454
rect 199794 489134 200414 489218
rect 199794 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 200414 489134
rect 199794 453454 200414 488898
rect 199794 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 200414 453454
rect 199794 453134 200414 453218
rect 199794 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 200414 453134
rect 199794 417454 200414 452898
rect 199794 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 200414 417454
rect 199794 417134 200414 417218
rect 199794 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 200414 417134
rect 199794 381454 200414 416898
rect 199794 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 200414 381454
rect 199794 381134 200414 381218
rect 199794 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 200414 381134
rect 199794 345454 200414 380898
rect 199794 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 200414 345454
rect 199794 345134 200414 345218
rect 199794 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 200414 345134
rect 199794 309454 200414 344898
rect 199794 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 200414 309454
rect 199794 309134 200414 309218
rect 199794 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 200414 309134
rect 199794 273454 200414 308898
rect 199794 273218 199826 273454
rect 200062 273218 200146 273454
rect 200382 273218 200414 273454
rect 199794 273134 200414 273218
rect 199794 272898 199826 273134
rect 200062 272898 200146 273134
rect 200382 272898 200414 273134
rect 199794 237454 200414 272898
rect 199794 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 200414 237454
rect 199794 237134 200414 237218
rect 199794 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 200414 237134
rect 199794 201454 200414 236898
rect 199794 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 200414 201454
rect 199794 201134 200414 201218
rect 199794 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 200414 201134
rect 199794 165454 200414 200898
rect 199794 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 200414 165454
rect 199794 165134 200414 165218
rect 199794 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 200414 165134
rect 199794 129454 200414 164898
rect 199794 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 200414 129454
rect 199794 129134 200414 129218
rect 199794 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 200414 129134
rect 199794 93454 200414 128898
rect 199794 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 200414 93454
rect 199794 93134 200414 93218
rect 199794 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 200414 93134
rect 199794 57454 200414 92898
rect 199794 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 200414 57454
rect 199794 57134 200414 57218
rect 199794 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 200414 57134
rect 199794 21454 200414 56898
rect 199794 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 200414 21454
rect 199794 21134 200414 21218
rect 199794 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 200414 21134
rect 199794 -4186 200414 20898
rect 199794 -4422 199826 -4186
rect 200062 -4422 200146 -4186
rect 200382 -4422 200414 -4186
rect 199794 -4506 200414 -4422
rect 199794 -4742 199826 -4506
rect 200062 -4742 200146 -4506
rect 200382 -4742 200414 -4506
rect 199794 -7654 200414 -4742
rect 204294 709638 204914 711590
rect 204294 709402 204326 709638
rect 204562 709402 204646 709638
rect 204882 709402 204914 709638
rect 204294 709318 204914 709402
rect 204294 709082 204326 709318
rect 204562 709082 204646 709318
rect 204882 709082 204914 709318
rect 204294 673954 204914 709082
rect 204294 673718 204326 673954
rect 204562 673718 204646 673954
rect 204882 673718 204914 673954
rect 204294 673634 204914 673718
rect 204294 673398 204326 673634
rect 204562 673398 204646 673634
rect 204882 673398 204914 673634
rect 204294 637954 204914 673398
rect 204294 637718 204326 637954
rect 204562 637718 204646 637954
rect 204882 637718 204914 637954
rect 204294 637634 204914 637718
rect 204294 637398 204326 637634
rect 204562 637398 204646 637634
rect 204882 637398 204914 637634
rect 204294 601954 204914 637398
rect 204294 601718 204326 601954
rect 204562 601718 204646 601954
rect 204882 601718 204914 601954
rect 204294 601634 204914 601718
rect 204294 601398 204326 601634
rect 204562 601398 204646 601634
rect 204882 601398 204914 601634
rect 204294 565954 204914 601398
rect 204294 565718 204326 565954
rect 204562 565718 204646 565954
rect 204882 565718 204914 565954
rect 204294 565634 204914 565718
rect 204294 565398 204326 565634
rect 204562 565398 204646 565634
rect 204882 565398 204914 565634
rect 204294 529954 204914 565398
rect 204294 529718 204326 529954
rect 204562 529718 204646 529954
rect 204882 529718 204914 529954
rect 204294 529634 204914 529718
rect 204294 529398 204326 529634
rect 204562 529398 204646 529634
rect 204882 529398 204914 529634
rect 204294 493954 204914 529398
rect 204294 493718 204326 493954
rect 204562 493718 204646 493954
rect 204882 493718 204914 493954
rect 204294 493634 204914 493718
rect 204294 493398 204326 493634
rect 204562 493398 204646 493634
rect 204882 493398 204914 493634
rect 204294 457954 204914 493398
rect 204294 457718 204326 457954
rect 204562 457718 204646 457954
rect 204882 457718 204914 457954
rect 204294 457634 204914 457718
rect 204294 457398 204326 457634
rect 204562 457398 204646 457634
rect 204882 457398 204914 457634
rect 204294 421954 204914 457398
rect 204294 421718 204326 421954
rect 204562 421718 204646 421954
rect 204882 421718 204914 421954
rect 204294 421634 204914 421718
rect 204294 421398 204326 421634
rect 204562 421398 204646 421634
rect 204882 421398 204914 421634
rect 204294 385954 204914 421398
rect 204294 385718 204326 385954
rect 204562 385718 204646 385954
rect 204882 385718 204914 385954
rect 204294 385634 204914 385718
rect 204294 385398 204326 385634
rect 204562 385398 204646 385634
rect 204882 385398 204914 385634
rect 204294 349954 204914 385398
rect 204294 349718 204326 349954
rect 204562 349718 204646 349954
rect 204882 349718 204914 349954
rect 204294 349634 204914 349718
rect 204294 349398 204326 349634
rect 204562 349398 204646 349634
rect 204882 349398 204914 349634
rect 204294 313954 204914 349398
rect 204294 313718 204326 313954
rect 204562 313718 204646 313954
rect 204882 313718 204914 313954
rect 204294 313634 204914 313718
rect 204294 313398 204326 313634
rect 204562 313398 204646 313634
rect 204882 313398 204914 313634
rect 204294 277954 204914 313398
rect 204294 277718 204326 277954
rect 204562 277718 204646 277954
rect 204882 277718 204914 277954
rect 204294 277634 204914 277718
rect 204294 277398 204326 277634
rect 204562 277398 204646 277634
rect 204882 277398 204914 277634
rect 204294 241954 204914 277398
rect 204294 241718 204326 241954
rect 204562 241718 204646 241954
rect 204882 241718 204914 241954
rect 204294 241634 204914 241718
rect 204294 241398 204326 241634
rect 204562 241398 204646 241634
rect 204882 241398 204914 241634
rect 204294 205954 204914 241398
rect 204294 205718 204326 205954
rect 204562 205718 204646 205954
rect 204882 205718 204914 205954
rect 204294 205634 204914 205718
rect 204294 205398 204326 205634
rect 204562 205398 204646 205634
rect 204882 205398 204914 205634
rect 204294 169954 204914 205398
rect 204294 169718 204326 169954
rect 204562 169718 204646 169954
rect 204882 169718 204914 169954
rect 204294 169634 204914 169718
rect 204294 169398 204326 169634
rect 204562 169398 204646 169634
rect 204882 169398 204914 169634
rect 204294 133954 204914 169398
rect 204294 133718 204326 133954
rect 204562 133718 204646 133954
rect 204882 133718 204914 133954
rect 204294 133634 204914 133718
rect 204294 133398 204326 133634
rect 204562 133398 204646 133634
rect 204882 133398 204914 133634
rect 204294 97954 204914 133398
rect 204294 97718 204326 97954
rect 204562 97718 204646 97954
rect 204882 97718 204914 97954
rect 204294 97634 204914 97718
rect 204294 97398 204326 97634
rect 204562 97398 204646 97634
rect 204882 97398 204914 97634
rect 204294 61954 204914 97398
rect 204294 61718 204326 61954
rect 204562 61718 204646 61954
rect 204882 61718 204914 61954
rect 204294 61634 204914 61718
rect 204294 61398 204326 61634
rect 204562 61398 204646 61634
rect 204882 61398 204914 61634
rect 204294 25954 204914 61398
rect 204294 25718 204326 25954
rect 204562 25718 204646 25954
rect 204882 25718 204914 25954
rect 204294 25634 204914 25718
rect 204294 25398 204326 25634
rect 204562 25398 204646 25634
rect 204882 25398 204914 25634
rect 204294 -5146 204914 25398
rect 204294 -5382 204326 -5146
rect 204562 -5382 204646 -5146
rect 204882 -5382 204914 -5146
rect 204294 -5466 204914 -5382
rect 204294 -5702 204326 -5466
rect 204562 -5702 204646 -5466
rect 204882 -5702 204914 -5466
rect 204294 -7654 204914 -5702
rect 208794 710598 209414 711590
rect 208794 710362 208826 710598
rect 209062 710362 209146 710598
rect 209382 710362 209414 710598
rect 208794 710278 209414 710362
rect 208794 710042 208826 710278
rect 209062 710042 209146 710278
rect 209382 710042 209414 710278
rect 208794 678454 209414 710042
rect 208794 678218 208826 678454
rect 209062 678218 209146 678454
rect 209382 678218 209414 678454
rect 208794 678134 209414 678218
rect 208794 677898 208826 678134
rect 209062 677898 209146 678134
rect 209382 677898 209414 678134
rect 208794 642454 209414 677898
rect 208794 642218 208826 642454
rect 209062 642218 209146 642454
rect 209382 642218 209414 642454
rect 208794 642134 209414 642218
rect 208794 641898 208826 642134
rect 209062 641898 209146 642134
rect 209382 641898 209414 642134
rect 208794 606454 209414 641898
rect 208794 606218 208826 606454
rect 209062 606218 209146 606454
rect 209382 606218 209414 606454
rect 208794 606134 209414 606218
rect 208794 605898 208826 606134
rect 209062 605898 209146 606134
rect 209382 605898 209414 606134
rect 208794 570454 209414 605898
rect 208794 570218 208826 570454
rect 209062 570218 209146 570454
rect 209382 570218 209414 570454
rect 208794 570134 209414 570218
rect 208794 569898 208826 570134
rect 209062 569898 209146 570134
rect 209382 569898 209414 570134
rect 208794 534454 209414 569898
rect 208794 534218 208826 534454
rect 209062 534218 209146 534454
rect 209382 534218 209414 534454
rect 208794 534134 209414 534218
rect 208794 533898 208826 534134
rect 209062 533898 209146 534134
rect 209382 533898 209414 534134
rect 208794 498454 209414 533898
rect 208794 498218 208826 498454
rect 209062 498218 209146 498454
rect 209382 498218 209414 498454
rect 208794 498134 209414 498218
rect 208794 497898 208826 498134
rect 209062 497898 209146 498134
rect 209382 497898 209414 498134
rect 208794 462454 209414 497898
rect 208794 462218 208826 462454
rect 209062 462218 209146 462454
rect 209382 462218 209414 462454
rect 208794 462134 209414 462218
rect 208794 461898 208826 462134
rect 209062 461898 209146 462134
rect 209382 461898 209414 462134
rect 208794 426454 209414 461898
rect 208794 426218 208826 426454
rect 209062 426218 209146 426454
rect 209382 426218 209414 426454
rect 208794 426134 209414 426218
rect 208794 425898 208826 426134
rect 209062 425898 209146 426134
rect 209382 425898 209414 426134
rect 208794 390454 209414 425898
rect 208794 390218 208826 390454
rect 209062 390218 209146 390454
rect 209382 390218 209414 390454
rect 208794 390134 209414 390218
rect 208794 389898 208826 390134
rect 209062 389898 209146 390134
rect 209382 389898 209414 390134
rect 208794 354454 209414 389898
rect 208794 354218 208826 354454
rect 209062 354218 209146 354454
rect 209382 354218 209414 354454
rect 208794 354134 209414 354218
rect 208794 353898 208826 354134
rect 209062 353898 209146 354134
rect 209382 353898 209414 354134
rect 208794 318454 209414 353898
rect 208794 318218 208826 318454
rect 209062 318218 209146 318454
rect 209382 318218 209414 318454
rect 208794 318134 209414 318218
rect 208794 317898 208826 318134
rect 209062 317898 209146 318134
rect 209382 317898 209414 318134
rect 208794 282454 209414 317898
rect 208794 282218 208826 282454
rect 209062 282218 209146 282454
rect 209382 282218 209414 282454
rect 208794 282134 209414 282218
rect 208794 281898 208826 282134
rect 209062 281898 209146 282134
rect 209382 281898 209414 282134
rect 208794 246454 209414 281898
rect 208794 246218 208826 246454
rect 209062 246218 209146 246454
rect 209382 246218 209414 246454
rect 208794 246134 209414 246218
rect 208794 245898 208826 246134
rect 209062 245898 209146 246134
rect 209382 245898 209414 246134
rect 208794 210454 209414 245898
rect 208794 210218 208826 210454
rect 209062 210218 209146 210454
rect 209382 210218 209414 210454
rect 208794 210134 209414 210218
rect 208794 209898 208826 210134
rect 209062 209898 209146 210134
rect 209382 209898 209414 210134
rect 208794 174454 209414 209898
rect 208794 174218 208826 174454
rect 209062 174218 209146 174454
rect 209382 174218 209414 174454
rect 208794 174134 209414 174218
rect 208794 173898 208826 174134
rect 209062 173898 209146 174134
rect 209382 173898 209414 174134
rect 208794 138454 209414 173898
rect 208794 138218 208826 138454
rect 209062 138218 209146 138454
rect 209382 138218 209414 138454
rect 208794 138134 209414 138218
rect 208794 137898 208826 138134
rect 209062 137898 209146 138134
rect 209382 137898 209414 138134
rect 208794 102454 209414 137898
rect 208794 102218 208826 102454
rect 209062 102218 209146 102454
rect 209382 102218 209414 102454
rect 208794 102134 209414 102218
rect 208794 101898 208826 102134
rect 209062 101898 209146 102134
rect 209382 101898 209414 102134
rect 208794 66454 209414 101898
rect 208794 66218 208826 66454
rect 209062 66218 209146 66454
rect 209382 66218 209414 66454
rect 208794 66134 209414 66218
rect 208794 65898 208826 66134
rect 209062 65898 209146 66134
rect 209382 65898 209414 66134
rect 208794 30454 209414 65898
rect 208794 30218 208826 30454
rect 209062 30218 209146 30454
rect 209382 30218 209414 30454
rect 208794 30134 209414 30218
rect 208794 29898 208826 30134
rect 209062 29898 209146 30134
rect 209382 29898 209414 30134
rect 208794 -6106 209414 29898
rect 208794 -6342 208826 -6106
rect 209062 -6342 209146 -6106
rect 209382 -6342 209414 -6106
rect 208794 -6426 209414 -6342
rect 208794 -6662 208826 -6426
rect 209062 -6662 209146 -6426
rect 209382 -6662 209414 -6426
rect 208794 -7654 209414 -6662
rect 213294 711558 213914 711590
rect 213294 711322 213326 711558
rect 213562 711322 213646 711558
rect 213882 711322 213914 711558
rect 213294 711238 213914 711322
rect 213294 711002 213326 711238
rect 213562 711002 213646 711238
rect 213882 711002 213914 711238
rect 213294 682954 213914 711002
rect 213294 682718 213326 682954
rect 213562 682718 213646 682954
rect 213882 682718 213914 682954
rect 213294 682634 213914 682718
rect 213294 682398 213326 682634
rect 213562 682398 213646 682634
rect 213882 682398 213914 682634
rect 213294 646954 213914 682398
rect 213294 646718 213326 646954
rect 213562 646718 213646 646954
rect 213882 646718 213914 646954
rect 213294 646634 213914 646718
rect 213294 646398 213326 646634
rect 213562 646398 213646 646634
rect 213882 646398 213914 646634
rect 213294 610954 213914 646398
rect 213294 610718 213326 610954
rect 213562 610718 213646 610954
rect 213882 610718 213914 610954
rect 213294 610634 213914 610718
rect 213294 610398 213326 610634
rect 213562 610398 213646 610634
rect 213882 610398 213914 610634
rect 213294 574954 213914 610398
rect 213294 574718 213326 574954
rect 213562 574718 213646 574954
rect 213882 574718 213914 574954
rect 213294 574634 213914 574718
rect 213294 574398 213326 574634
rect 213562 574398 213646 574634
rect 213882 574398 213914 574634
rect 213294 538954 213914 574398
rect 213294 538718 213326 538954
rect 213562 538718 213646 538954
rect 213882 538718 213914 538954
rect 213294 538634 213914 538718
rect 213294 538398 213326 538634
rect 213562 538398 213646 538634
rect 213882 538398 213914 538634
rect 213294 502954 213914 538398
rect 213294 502718 213326 502954
rect 213562 502718 213646 502954
rect 213882 502718 213914 502954
rect 213294 502634 213914 502718
rect 213294 502398 213326 502634
rect 213562 502398 213646 502634
rect 213882 502398 213914 502634
rect 213294 466954 213914 502398
rect 213294 466718 213326 466954
rect 213562 466718 213646 466954
rect 213882 466718 213914 466954
rect 213294 466634 213914 466718
rect 213294 466398 213326 466634
rect 213562 466398 213646 466634
rect 213882 466398 213914 466634
rect 213294 430954 213914 466398
rect 213294 430718 213326 430954
rect 213562 430718 213646 430954
rect 213882 430718 213914 430954
rect 213294 430634 213914 430718
rect 213294 430398 213326 430634
rect 213562 430398 213646 430634
rect 213882 430398 213914 430634
rect 213294 394954 213914 430398
rect 213294 394718 213326 394954
rect 213562 394718 213646 394954
rect 213882 394718 213914 394954
rect 213294 394634 213914 394718
rect 213294 394398 213326 394634
rect 213562 394398 213646 394634
rect 213882 394398 213914 394634
rect 213294 358954 213914 394398
rect 213294 358718 213326 358954
rect 213562 358718 213646 358954
rect 213882 358718 213914 358954
rect 213294 358634 213914 358718
rect 213294 358398 213326 358634
rect 213562 358398 213646 358634
rect 213882 358398 213914 358634
rect 213294 322954 213914 358398
rect 213294 322718 213326 322954
rect 213562 322718 213646 322954
rect 213882 322718 213914 322954
rect 213294 322634 213914 322718
rect 213294 322398 213326 322634
rect 213562 322398 213646 322634
rect 213882 322398 213914 322634
rect 213294 286954 213914 322398
rect 213294 286718 213326 286954
rect 213562 286718 213646 286954
rect 213882 286718 213914 286954
rect 213294 286634 213914 286718
rect 213294 286398 213326 286634
rect 213562 286398 213646 286634
rect 213882 286398 213914 286634
rect 213294 250954 213914 286398
rect 213294 250718 213326 250954
rect 213562 250718 213646 250954
rect 213882 250718 213914 250954
rect 213294 250634 213914 250718
rect 213294 250398 213326 250634
rect 213562 250398 213646 250634
rect 213882 250398 213914 250634
rect 213294 214954 213914 250398
rect 213294 214718 213326 214954
rect 213562 214718 213646 214954
rect 213882 214718 213914 214954
rect 213294 214634 213914 214718
rect 213294 214398 213326 214634
rect 213562 214398 213646 214634
rect 213882 214398 213914 214634
rect 213294 178954 213914 214398
rect 213294 178718 213326 178954
rect 213562 178718 213646 178954
rect 213882 178718 213914 178954
rect 213294 178634 213914 178718
rect 213294 178398 213326 178634
rect 213562 178398 213646 178634
rect 213882 178398 213914 178634
rect 213294 142954 213914 178398
rect 213294 142718 213326 142954
rect 213562 142718 213646 142954
rect 213882 142718 213914 142954
rect 213294 142634 213914 142718
rect 213294 142398 213326 142634
rect 213562 142398 213646 142634
rect 213882 142398 213914 142634
rect 213294 106954 213914 142398
rect 213294 106718 213326 106954
rect 213562 106718 213646 106954
rect 213882 106718 213914 106954
rect 213294 106634 213914 106718
rect 213294 106398 213326 106634
rect 213562 106398 213646 106634
rect 213882 106398 213914 106634
rect 213294 70954 213914 106398
rect 213294 70718 213326 70954
rect 213562 70718 213646 70954
rect 213882 70718 213914 70954
rect 213294 70634 213914 70718
rect 213294 70398 213326 70634
rect 213562 70398 213646 70634
rect 213882 70398 213914 70634
rect 213294 34954 213914 70398
rect 213294 34718 213326 34954
rect 213562 34718 213646 34954
rect 213882 34718 213914 34954
rect 213294 34634 213914 34718
rect 213294 34398 213326 34634
rect 213562 34398 213646 34634
rect 213882 34398 213914 34634
rect 213294 -7066 213914 34398
rect 213294 -7302 213326 -7066
rect 213562 -7302 213646 -7066
rect 213882 -7302 213914 -7066
rect 213294 -7386 213914 -7302
rect 213294 -7622 213326 -7386
rect 213562 -7622 213646 -7386
rect 213882 -7622 213914 -7386
rect 213294 -7654 213914 -7622
rect 217794 704838 218414 711590
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 687454 218414 704282
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 651454 218414 686898
rect 217794 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 218414 651454
rect 217794 651134 218414 651218
rect 217794 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 218414 651134
rect 217794 615454 218414 650898
rect 217794 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 218414 615454
rect 217794 615134 218414 615218
rect 217794 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 218414 615134
rect 217794 579454 218414 614898
rect 217794 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 218414 579454
rect 217794 579134 218414 579218
rect 217794 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 218414 579134
rect 217794 543454 218414 578898
rect 217794 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 218414 543454
rect 217794 543134 218414 543218
rect 217794 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 218414 543134
rect 217794 507454 218414 542898
rect 217794 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 218414 507454
rect 217794 507134 218414 507218
rect 217794 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 218414 507134
rect 217794 471454 218414 506898
rect 217794 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 218414 471454
rect 217794 471134 218414 471218
rect 217794 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 218414 471134
rect 217794 435454 218414 470898
rect 217794 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 218414 435454
rect 217794 435134 218414 435218
rect 217794 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 218414 435134
rect 217794 399454 218414 434898
rect 217794 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 218414 399454
rect 217794 399134 218414 399218
rect 217794 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 218414 399134
rect 217794 363454 218414 398898
rect 217794 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 218414 363454
rect 217794 363134 218414 363218
rect 217794 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 218414 363134
rect 217794 327454 218414 362898
rect 217794 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 218414 327454
rect 217794 327134 218414 327218
rect 217794 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 218414 327134
rect 217794 291454 218414 326898
rect 217794 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 218414 291454
rect 217794 291134 218414 291218
rect 217794 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 218414 291134
rect 217794 255454 218414 290898
rect 217794 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 218414 255454
rect 217794 255134 218414 255218
rect 217794 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 218414 255134
rect 217794 219454 218414 254898
rect 217794 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 218414 219454
rect 217794 219134 218414 219218
rect 217794 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 218414 219134
rect 217794 183454 218414 218898
rect 217794 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 218414 183454
rect 217794 183134 218414 183218
rect 217794 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 218414 183134
rect 217794 147454 218414 182898
rect 217794 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 218414 147454
rect 217794 147134 218414 147218
rect 217794 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 218414 147134
rect 217794 111454 218414 146898
rect 217794 111218 217826 111454
rect 218062 111218 218146 111454
rect 218382 111218 218414 111454
rect 217794 111134 218414 111218
rect 217794 110898 217826 111134
rect 218062 110898 218146 111134
rect 218382 110898 218414 111134
rect 217794 75454 218414 110898
rect 217794 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 218414 75454
rect 217794 75134 218414 75218
rect 217794 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 218414 75134
rect 217794 39454 218414 74898
rect 217794 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 218414 39454
rect 217794 39134 218414 39218
rect 217794 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 218414 39134
rect 217794 3454 218414 38898
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -7654 218414 -902
rect 222294 705798 222914 711590
rect 222294 705562 222326 705798
rect 222562 705562 222646 705798
rect 222882 705562 222914 705798
rect 222294 705478 222914 705562
rect 222294 705242 222326 705478
rect 222562 705242 222646 705478
rect 222882 705242 222914 705478
rect 222294 691954 222914 705242
rect 222294 691718 222326 691954
rect 222562 691718 222646 691954
rect 222882 691718 222914 691954
rect 222294 691634 222914 691718
rect 222294 691398 222326 691634
rect 222562 691398 222646 691634
rect 222882 691398 222914 691634
rect 222294 655954 222914 691398
rect 222294 655718 222326 655954
rect 222562 655718 222646 655954
rect 222882 655718 222914 655954
rect 222294 655634 222914 655718
rect 222294 655398 222326 655634
rect 222562 655398 222646 655634
rect 222882 655398 222914 655634
rect 222294 619954 222914 655398
rect 222294 619718 222326 619954
rect 222562 619718 222646 619954
rect 222882 619718 222914 619954
rect 222294 619634 222914 619718
rect 222294 619398 222326 619634
rect 222562 619398 222646 619634
rect 222882 619398 222914 619634
rect 222294 583954 222914 619398
rect 222294 583718 222326 583954
rect 222562 583718 222646 583954
rect 222882 583718 222914 583954
rect 222294 583634 222914 583718
rect 222294 583398 222326 583634
rect 222562 583398 222646 583634
rect 222882 583398 222914 583634
rect 222294 547954 222914 583398
rect 222294 547718 222326 547954
rect 222562 547718 222646 547954
rect 222882 547718 222914 547954
rect 222294 547634 222914 547718
rect 222294 547398 222326 547634
rect 222562 547398 222646 547634
rect 222882 547398 222914 547634
rect 222294 511954 222914 547398
rect 222294 511718 222326 511954
rect 222562 511718 222646 511954
rect 222882 511718 222914 511954
rect 222294 511634 222914 511718
rect 222294 511398 222326 511634
rect 222562 511398 222646 511634
rect 222882 511398 222914 511634
rect 222294 475954 222914 511398
rect 222294 475718 222326 475954
rect 222562 475718 222646 475954
rect 222882 475718 222914 475954
rect 222294 475634 222914 475718
rect 222294 475398 222326 475634
rect 222562 475398 222646 475634
rect 222882 475398 222914 475634
rect 222294 439954 222914 475398
rect 222294 439718 222326 439954
rect 222562 439718 222646 439954
rect 222882 439718 222914 439954
rect 222294 439634 222914 439718
rect 222294 439398 222326 439634
rect 222562 439398 222646 439634
rect 222882 439398 222914 439634
rect 222294 403954 222914 439398
rect 222294 403718 222326 403954
rect 222562 403718 222646 403954
rect 222882 403718 222914 403954
rect 222294 403634 222914 403718
rect 222294 403398 222326 403634
rect 222562 403398 222646 403634
rect 222882 403398 222914 403634
rect 222294 367954 222914 403398
rect 222294 367718 222326 367954
rect 222562 367718 222646 367954
rect 222882 367718 222914 367954
rect 222294 367634 222914 367718
rect 222294 367398 222326 367634
rect 222562 367398 222646 367634
rect 222882 367398 222914 367634
rect 222294 331954 222914 367398
rect 222294 331718 222326 331954
rect 222562 331718 222646 331954
rect 222882 331718 222914 331954
rect 222294 331634 222914 331718
rect 222294 331398 222326 331634
rect 222562 331398 222646 331634
rect 222882 331398 222914 331634
rect 222294 295954 222914 331398
rect 222294 295718 222326 295954
rect 222562 295718 222646 295954
rect 222882 295718 222914 295954
rect 222294 295634 222914 295718
rect 222294 295398 222326 295634
rect 222562 295398 222646 295634
rect 222882 295398 222914 295634
rect 222294 259954 222914 295398
rect 222294 259718 222326 259954
rect 222562 259718 222646 259954
rect 222882 259718 222914 259954
rect 222294 259634 222914 259718
rect 222294 259398 222326 259634
rect 222562 259398 222646 259634
rect 222882 259398 222914 259634
rect 222294 223954 222914 259398
rect 222294 223718 222326 223954
rect 222562 223718 222646 223954
rect 222882 223718 222914 223954
rect 222294 223634 222914 223718
rect 222294 223398 222326 223634
rect 222562 223398 222646 223634
rect 222882 223398 222914 223634
rect 222294 187954 222914 223398
rect 222294 187718 222326 187954
rect 222562 187718 222646 187954
rect 222882 187718 222914 187954
rect 222294 187634 222914 187718
rect 222294 187398 222326 187634
rect 222562 187398 222646 187634
rect 222882 187398 222914 187634
rect 222294 151954 222914 187398
rect 222294 151718 222326 151954
rect 222562 151718 222646 151954
rect 222882 151718 222914 151954
rect 222294 151634 222914 151718
rect 222294 151398 222326 151634
rect 222562 151398 222646 151634
rect 222882 151398 222914 151634
rect 222294 115954 222914 151398
rect 222294 115718 222326 115954
rect 222562 115718 222646 115954
rect 222882 115718 222914 115954
rect 222294 115634 222914 115718
rect 222294 115398 222326 115634
rect 222562 115398 222646 115634
rect 222882 115398 222914 115634
rect 222294 79954 222914 115398
rect 222294 79718 222326 79954
rect 222562 79718 222646 79954
rect 222882 79718 222914 79954
rect 222294 79634 222914 79718
rect 222294 79398 222326 79634
rect 222562 79398 222646 79634
rect 222882 79398 222914 79634
rect 222294 43954 222914 79398
rect 222294 43718 222326 43954
rect 222562 43718 222646 43954
rect 222882 43718 222914 43954
rect 222294 43634 222914 43718
rect 222294 43398 222326 43634
rect 222562 43398 222646 43634
rect 222882 43398 222914 43634
rect 222294 7954 222914 43398
rect 222294 7718 222326 7954
rect 222562 7718 222646 7954
rect 222882 7718 222914 7954
rect 222294 7634 222914 7718
rect 222294 7398 222326 7634
rect 222562 7398 222646 7634
rect 222882 7398 222914 7634
rect 222294 -1306 222914 7398
rect 222294 -1542 222326 -1306
rect 222562 -1542 222646 -1306
rect 222882 -1542 222914 -1306
rect 222294 -1626 222914 -1542
rect 222294 -1862 222326 -1626
rect 222562 -1862 222646 -1626
rect 222882 -1862 222914 -1626
rect 222294 -7654 222914 -1862
rect 226794 706758 227414 711590
rect 226794 706522 226826 706758
rect 227062 706522 227146 706758
rect 227382 706522 227414 706758
rect 226794 706438 227414 706522
rect 226794 706202 226826 706438
rect 227062 706202 227146 706438
rect 227382 706202 227414 706438
rect 226794 696454 227414 706202
rect 226794 696218 226826 696454
rect 227062 696218 227146 696454
rect 227382 696218 227414 696454
rect 226794 696134 227414 696218
rect 226794 695898 226826 696134
rect 227062 695898 227146 696134
rect 227382 695898 227414 696134
rect 226794 660454 227414 695898
rect 226794 660218 226826 660454
rect 227062 660218 227146 660454
rect 227382 660218 227414 660454
rect 226794 660134 227414 660218
rect 226794 659898 226826 660134
rect 227062 659898 227146 660134
rect 227382 659898 227414 660134
rect 226794 624454 227414 659898
rect 226794 624218 226826 624454
rect 227062 624218 227146 624454
rect 227382 624218 227414 624454
rect 226794 624134 227414 624218
rect 226794 623898 226826 624134
rect 227062 623898 227146 624134
rect 227382 623898 227414 624134
rect 226794 588454 227414 623898
rect 226794 588218 226826 588454
rect 227062 588218 227146 588454
rect 227382 588218 227414 588454
rect 226794 588134 227414 588218
rect 226794 587898 226826 588134
rect 227062 587898 227146 588134
rect 227382 587898 227414 588134
rect 226794 552454 227414 587898
rect 226794 552218 226826 552454
rect 227062 552218 227146 552454
rect 227382 552218 227414 552454
rect 226794 552134 227414 552218
rect 226794 551898 226826 552134
rect 227062 551898 227146 552134
rect 227382 551898 227414 552134
rect 226794 516454 227414 551898
rect 226794 516218 226826 516454
rect 227062 516218 227146 516454
rect 227382 516218 227414 516454
rect 226794 516134 227414 516218
rect 226794 515898 226826 516134
rect 227062 515898 227146 516134
rect 227382 515898 227414 516134
rect 226794 480454 227414 515898
rect 226794 480218 226826 480454
rect 227062 480218 227146 480454
rect 227382 480218 227414 480454
rect 226794 480134 227414 480218
rect 226794 479898 226826 480134
rect 227062 479898 227146 480134
rect 227382 479898 227414 480134
rect 226794 444454 227414 479898
rect 226794 444218 226826 444454
rect 227062 444218 227146 444454
rect 227382 444218 227414 444454
rect 226794 444134 227414 444218
rect 226794 443898 226826 444134
rect 227062 443898 227146 444134
rect 227382 443898 227414 444134
rect 226794 408454 227414 443898
rect 226794 408218 226826 408454
rect 227062 408218 227146 408454
rect 227382 408218 227414 408454
rect 226794 408134 227414 408218
rect 226794 407898 226826 408134
rect 227062 407898 227146 408134
rect 227382 407898 227414 408134
rect 226794 372454 227414 407898
rect 226794 372218 226826 372454
rect 227062 372218 227146 372454
rect 227382 372218 227414 372454
rect 226794 372134 227414 372218
rect 226794 371898 226826 372134
rect 227062 371898 227146 372134
rect 227382 371898 227414 372134
rect 226794 336454 227414 371898
rect 226794 336218 226826 336454
rect 227062 336218 227146 336454
rect 227382 336218 227414 336454
rect 226794 336134 227414 336218
rect 226794 335898 226826 336134
rect 227062 335898 227146 336134
rect 227382 335898 227414 336134
rect 226794 300454 227414 335898
rect 226794 300218 226826 300454
rect 227062 300218 227146 300454
rect 227382 300218 227414 300454
rect 226794 300134 227414 300218
rect 226794 299898 226826 300134
rect 227062 299898 227146 300134
rect 227382 299898 227414 300134
rect 226794 264454 227414 299898
rect 226794 264218 226826 264454
rect 227062 264218 227146 264454
rect 227382 264218 227414 264454
rect 226794 264134 227414 264218
rect 226794 263898 226826 264134
rect 227062 263898 227146 264134
rect 227382 263898 227414 264134
rect 226794 228454 227414 263898
rect 226794 228218 226826 228454
rect 227062 228218 227146 228454
rect 227382 228218 227414 228454
rect 226794 228134 227414 228218
rect 226794 227898 226826 228134
rect 227062 227898 227146 228134
rect 227382 227898 227414 228134
rect 226794 192454 227414 227898
rect 226794 192218 226826 192454
rect 227062 192218 227146 192454
rect 227382 192218 227414 192454
rect 226794 192134 227414 192218
rect 226794 191898 226826 192134
rect 227062 191898 227146 192134
rect 227382 191898 227414 192134
rect 226794 156454 227414 191898
rect 226794 156218 226826 156454
rect 227062 156218 227146 156454
rect 227382 156218 227414 156454
rect 226794 156134 227414 156218
rect 226794 155898 226826 156134
rect 227062 155898 227146 156134
rect 227382 155898 227414 156134
rect 226794 120454 227414 155898
rect 226794 120218 226826 120454
rect 227062 120218 227146 120454
rect 227382 120218 227414 120454
rect 226794 120134 227414 120218
rect 226794 119898 226826 120134
rect 227062 119898 227146 120134
rect 227382 119898 227414 120134
rect 226794 84454 227414 119898
rect 226794 84218 226826 84454
rect 227062 84218 227146 84454
rect 227382 84218 227414 84454
rect 226794 84134 227414 84218
rect 226794 83898 226826 84134
rect 227062 83898 227146 84134
rect 227382 83898 227414 84134
rect 226794 48454 227414 83898
rect 226794 48218 226826 48454
rect 227062 48218 227146 48454
rect 227382 48218 227414 48454
rect 226794 48134 227414 48218
rect 226794 47898 226826 48134
rect 227062 47898 227146 48134
rect 227382 47898 227414 48134
rect 226794 12454 227414 47898
rect 226794 12218 226826 12454
rect 227062 12218 227146 12454
rect 227382 12218 227414 12454
rect 226794 12134 227414 12218
rect 226794 11898 226826 12134
rect 227062 11898 227146 12134
rect 227382 11898 227414 12134
rect 226794 -2266 227414 11898
rect 226794 -2502 226826 -2266
rect 227062 -2502 227146 -2266
rect 227382 -2502 227414 -2266
rect 226794 -2586 227414 -2502
rect 226794 -2822 226826 -2586
rect 227062 -2822 227146 -2586
rect 227382 -2822 227414 -2586
rect 226794 -7654 227414 -2822
rect 231294 707718 231914 711590
rect 231294 707482 231326 707718
rect 231562 707482 231646 707718
rect 231882 707482 231914 707718
rect 231294 707398 231914 707482
rect 231294 707162 231326 707398
rect 231562 707162 231646 707398
rect 231882 707162 231914 707398
rect 231294 700954 231914 707162
rect 231294 700718 231326 700954
rect 231562 700718 231646 700954
rect 231882 700718 231914 700954
rect 231294 700634 231914 700718
rect 231294 700398 231326 700634
rect 231562 700398 231646 700634
rect 231882 700398 231914 700634
rect 231294 664954 231914 700398
rect 231294 664718 231326 664954
rect 231562 664718 231646 664954
rect 231882 664718 231914 664954
rect 231294 664634 231914 664718
rect 231294 664398 231326 664634
rect 231562 664398 231646 664634
rect 231882 664398 231914 664634
rect 231294 628954 231914 664398
rect 231294 628718 231326 628954
rect 231562 628718 231646 628954
rect 231882 628718 231914 628954
rect 231294 628634 231914 628718
rect 231294 628398 231326 628634
rect 231562 628398 231646 628634
rect 231882 628398 231914 628634
rect 231294 592954 231914 628398
rect 231294 592718 231326 592954
rect 231562 592718 231646 592954
rect 231882 592718 231914 592954
rect 231294 592634 231914 592718
rect 231294 592398 231326 592634
rect 231562 592398 231646 592634
rect 231882 592398 231914 592634
rect 231294 556954 231914 592398
rect 231294 556718 231326 556954
rect 231562 556718 231646 556954
rect 231882 556718 231914 556954
rect 231294 556634 231914 556718
rect 231294 556398 231326 556634
rect 231562 556398 231646 556634
rect 231882 556398 231914 556634
rect 231294 520954 231914 556398
rect 231294 520718 231326 520954
rect 231562 520718 231646 520954
rect 231882 520718 231914 520954
rect 231294 520634 231914 520718
rect 231294 520398 231326 520634
rect 231562 520398 231646 520634
rect 231882 520398 231914 520634
rect 231294 484954 231914 520398
rect 231294 484718 231326 484954
rect 231562 484718 231646 484954
rect 231882 484718 231914 484954
rect 231294 484634 231914 484718
rect 231294 484398 231326 484634
rect 231562 484398 231646 484634
rect 231882 484398 231914 484634
rect 231294 448954 231914 484398
rect 231294 448718 231326 448954
rect 231562 448718 231646 448954
rect 231882 448718 231914 448954
rect 231294 448634 231914 448718
rect 231294 448398 231326 448634
rect 231562 448398 231646 448634
rect 231882 448398 231914 448634
rect 231294 412954 231914 448398
rect 231294 412718 231326 412954
rect 231562 412718 231646 412954
rect 231882 412718 231914 412954
rect 231294 412634 231914 412718
rect 231294 412398 231326 412634
rect 231562 412398 231646 412634
rect 231882 412398 231914 412634
rect 231294 376954 231914 412398
rect 235794 708678 236414 711590
rect 235794 708442 235826 708678
rect 236062 708442 236146 708678
rect 236382 708442 236414 708678
rect 235794 708358 236414 708442
rect 235794 708122 235826 708358
rect 236062 708122 236146 708358
rect 236382 708122 236414 708358
rect 235794 669454 236414 708122
rect 235794 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 236414 669454
rect 235794 669134 236414 669218
rect 235794 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 236414 669134
rect 235794 633454 236414 668898
rect 235794 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 236414 633454
rect 235794 633134 236414 633218
rect 235794 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 236414 633134
rect 235794 597454 236414 632898
rect 235794 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 236414 597454
rect 235794 597134 236414 597218
rect 235794 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 236414 597134
rect 235794 561454 236414 596898
rect 235794 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 236414 561454
rect 235794 561134 236414 561218
rect 235794 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 236414 561134
rect 235794 525454 236414 560898
rect 235794 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 236414 525454
rect 235794 525134 236414 525218
rect 235794 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 236414 525134
rect 235794 489454 236414 524898
rect 235794 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 236414 489454
rect 235794 489134 236414 489218
rect 235794 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 236414 489134
rect 235794 453454 236414 488898
rect 235794 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 236414 453454
rect 235794 453134 236414 453218
rect 235794 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 236414 453134
rect 235794 417454 236414 452898
rect 235794 417218 235826 417454
rect 236062 417218 236146 417454
rect 236382 417218 236414 417454
rect 235794 417134 236414 417218
rect 235794 416898 235826 417134
rect 236062 416898 236146 417134
rect 236382 416898 236414 417134
rect 233739 393412 233805 393413
rect 233739 393348 233740 393412
rect 233804 393348 233805 393412
rect 233739 393347 233805 393348
rect 231294 376718 231326 376954
rect 231562 376718 231646 376954
rect 231882 376718 231914 376954
rect 231294 376634 231914 376718
rect 231294 376398 231326 376634
rect 231562 376398 231646 376634
rect 231882 376398 231914 376634
rect 231294 340954 231914 376398
rect 231294 340718 231326 340954
rect 231562 340718 231646 340954
rect 231882 340718 231914 340954
rect 231294 340634 231914 340718
rect 231294 340398 231326 340634
rect 231562 340398 231646 340634
rect 231882 340398 231914 340634
rect 231294 304954 231914 340398
rect 231294 304718 231326 304954
rect 231562 304718 231646 304954
rect 231882 304718 231914 304954
rect 231294 304634 231914 304718
rect 231294 304398 231326 304634
rect 231562 304398 231646 304634
rect 231882 304398 231914 304634
rect 231294 268954 231914 304398
rect 231294 268718 231326 268954
rect 231562 268718 231646 268954
rect 231882 268718 231914 268954
rect 231294 268634 231914 268718
rect 231294 268398 231326 268634
rect 231562 268398 231646 268634
rect 231882 268398 231914 268634
rect 231294 232954 231914 268398
rect 231294 232718 231326 232954
rect 231562 232718 231646 232954
rect 231882 232718 231914 232954
rect 231294 232634 231914 232718
rect 231294 232398 231326 232634
rect 231562 232398 231646 232634
rect 231882 232398 231914 232634
rect 231294 196954 231914 232398
rect 231294 196718 231326 196954
rect 231562 196718 231646 196954
rect 231882 196718 231914 196954
rect 231294 196634 231914 196718
rect 231294 196398 231326 196634
rect 231562 196398 231646 196634
rect 231882 196398 231914 196634
rect 231294 160954 231914 196398
rect 231294 160718 231326 160954
rect 231562 160718 231646 160954
rect 231882 160718 231914 160954
rect 231294 160634 231914 160718
rect 231294 160398 231326 160634
rect 231562 160398 231646 160634
rect 231882 160398 231914 160634
rect 231294 124954 231914 160398
rect 231294 124718 231326 124954
rect 231562 124718 231646 124954
rect 231882 124718 231914 124954
rect 231294 124634 231914 124718
rect 231294 124398 231326 124634
rect 231562 124398 231646 124634
rect 231882 124398 231914 124634
rect 231294 88954 231914 124398
rect 233742 97885 233802 393347
rect 235211 384028 235277 384029
rect 235211 383964 235212 384028
rect 235276 383964 235277 384028
rect 235794 384000 236414 416898
rect 240294 709638 240914 711590
rect 240294 709402 240326 709638
rect 240562 709402 240646 709638
rect 240882 709402 240914 709638
rect 240294 709318 240914 709402
rect 240294 709082 240326 709318
rect 240562 709082 240646 709318
rect 240882 709082 240914 709318
rect 240294 673954 240914 709082
rect 240294 673718 240326 673954
rect 240562 673718 240646 673954
rect 240882 673718 240914 673954
rect 240294 673634 240914 673718
rect 240294 673398 240326 673634
rect 240562 673398 240646 673634
rect 240882 673398 240914 673634
rect 240294 637954 240914 673398
rect 240294 637718 240326 637954
rect 240562 637718 240646 637954
rect 240882 637718 240914 637954
rect 240294 637634 240914 637718
rect 240294 637398 240326 637634
rect 240562 637398 240646 637634
rect 240882 637398 240914 637634
rect 240294 601954 240914 637398
rect 240294 601718 240326 601954
rect 240562 601718 240646 601954
rect 240882 601718 240914 601954
rect 240294 601634 240914 601718
rect 240294 601398 240326 601634
rect 240562 601398 240646 601634
rect 240882 601398 240914 601634
rect 240294 565954 240914 601398
rect 240294 565718 240326 565954
rect 240562 565718 240646 565954
rect 240882 565718 240914 565954
rect 240294 565634 240914 565718
rect 240294 565398 240326 565634
rect 240562 565398 240646 565634
rect 240882 565398 240914 565634
rect 240294 529954 240914 565398
rect 240294 529718 240326 529954
rect 240562 529718 240646 529954
rect 240882 529718 240914 529954
rect 240294 529634 240914 529718
rect 240294 529398 240326 529634
rect 240562 529398 240646 529634
rect 240882 529398 240914 529634
rect 240294 493954 240914 529398
rect 240294 493718 240326 493954
rect 240562 493718 240646 493954
rect 240882 493718 240914 493954
rect 240294 493634 240914 493718
rect 240294 493398 240326 493634
rect 240562 493398 240646 493634
rect 240882 493398 240914 493634
rect 240294 457954 240914 493398
rect 240294 457718 240326 457954
rect 240562 457718 240646 457954
rect 240882 457718 240914 457954
rect 240294 457634 240914 457718
rect 240294 457398 240326 457634
rect 240562 457398 240646 457634
rect 240882 457398 240914 457634
rect 240294 421954 240914 457398
rect 240294 421718 240326 421954
rect 240562 421718 240646 421954
rect 240882 421718 240914 421954
rect 240294 421634 240914 421718
rect 240294 421398 240326 421634
rect 240562 421398 240646 421634
rect 240882 421398 240914 421634
rect 240294 385954 240914 421398
rect 240294 385718 240326 385954
rect 240562 385718 240646 385954
rect 240882 385718 240914 385954
rect 240294 385634 240914 385718
rect 240294 385398 240326 385634
rect 240562 385398 240646 385634
rect 240882 385398 240914 385634
rect 239627 385116 239693 385117
rect 239627 385052 239628 385116
rect 239692 385052 239693 385116
rect 239627 385051 239693 385052
rect 238523 384572 238589 384573
rect 238523 384508 238524 384572
rect 238588 384508 238589 384572
rect 238523 384507 238589 384508
rect 238155 384164 238221 384165
rect 238155 384100 238156 384164
rect 238220 384100 238221 384164
rect 238155 384099 238221 384100
rect 235211 383963 235277 383964
rect 233739 97884 233805 97885
rect 233739 97820 233740 97884
rect 233804 97820 233805 97884
rect 233739 97819 233805 97820
rect 235214 96661 235274 383963
rect 237235 381852 237301 381853
rect 237235 381788 237236 381852
rect 237300 381788 237301 381852
rect 237235 381787 237301 381788
rect 237051 380628 237117 380629
rect 237051 380564 237052 380628
rect 237116 380564 237117 380628
rect 237051 380563 237117 380564
rect 235794 309454 236414 336000
rect 235794 309218 235826 309454
rect 236062 309218 236146 309454
rect 236382 309218 236414 309454
rect 235794 309134 236414 309218
rect 235794 308898 235826 309134
rect 236062 308898 236146 309134
rect 236382 308898 236414 309134
rect 235794 273454 236414 308898
rect 235794 273218 235826 273454
rect 236062 273218 236146 273454
rect 236382 273218 236414 273454
rect 235794 273134 236414 273218
rect 235794 272898 235826 273134
rect 236062 272898 236146 273134
rect 236382 272898 236414 273134
rect 235794 237454 236414 272898
rect 235794 237218 235826 237454
rect 236062 237218 236146 237454
rect 236382 237218 236414 237454
rect 235794 237134 236414 237218
rect 235794 236898 235826 237134
rect 236062 236898 236146 237134
rect 236382 236898 236414 237134
rect 235794 201454 236414 236898
rect 235794 201218 235826 201454
rect 236062 201218 236146 201454
rect 236382 201218 236414 201454
rect 235794 201134 236414 201218
rect 235794 200898 235826 201134
rect 236062 200898 236146 201134
rect 236382 200898 236414 201134
rect 235794 165454 236414 200898
rect 235794 165218 235826 165454
rect 236062 165218 236146 165454
rect 236382 165218 236414 165454
rect 235794 165134 236414 165218
rect 235794 164898 235826 165134
rect 236062 164898 236146 165134
rect 236382 164898 236414 165134
rect 235794 129454 236414 164898
rect 235794 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 236414 129454
rect 235794 129134 236414 129218
rect 235794 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 236414 129134
rect 235211 96660 235277 96661
rect 235211 96596 235212 96660
rect 235276 96596 235277 96660
rect 235211 96595 235277 96596
rect 231294 88718 231326 88954
rect 231562 88718 231646 88954
rect 231882 88718 231914 88954
rect 231294 88634 231914 88718
rect 231294 88398 231326 88634
rect 231562 88398 231646 88634
rect 231882 88398 231914 88634
rect 231294 52954 231914 88398
rect 231294 52718 231326 52954
rect 231562 52718 231646 52954
rect 231882 52718 231914 52954
rect 231294 52634 231914 52718
rect 231294 52398 231326 52634
rect 231562 52398 231646 52634
rect 231882 52398 231914 52634
rect 231294 16954 231914 52398
rect 231294 16718 231326 16954
rect 231562 16718 231646 16954
rect 231882 16718 231914 16954
rect 231294 16634 231914 16718
rect 231294 16398 231326 16634
rect 231562 16398 231646 16634
rect 231882 16398 231914 16634
rect 231294 -3226 231914 16398
rect 231294 -3462 231326 -3226
rect 231562 -3462 231646 -3226
rect 231882 -3462 231914 -3226
rect 231294 -3546 231914 -3462
rect 231294 -3782 231326 -3546
rect 231562 -3782 231646 -3546
rect 231882 -3782 231914 -3546
rect 231294 -7654 231914 -3782
rect 235794 93454 236414 128898
rect 237054 115973 237114 380563
rect 237051 115972 237117 115973
rect 237051 115908 237052 115972
rect 237116 115908 237117 115972
rect 237051 115907 237117 115908
rect 237238 97613 237298 381787
rect 238158 214573 238218 384099
rect 238339 363492 238405 363493
rect 238339 363428 238340 363492
rect 238404 363428 238405 363492
rect 238339 363427 238405 363428
rect 238155 214572 238221 214573
rect 238155 214508 238156 214572
rect 238220 214508 238221 214572
rect 238155 214507 238221 214508
rect 238342 97749 238402 363427
rect 238526 107677 238586 384507
rect 238891 363492 238957 363493
rect 238891 363428 238892 363492
rect 238956 363428 238957 363492
rect 238891 363427 238957 363428
rect 239208 363454 239528 363486
rect 238894 339965 238954 363427
rect 239208 363218 239250 363454
rect 239486 363218 239528 363454
rect 239208 363134 239528 363218
rect 239208 362898 239250 363134
rect 239486 362898 239528 363134
rect 239208 362866 239528 362898
rect 239630 339965 239690 385051
rect 240294 384000 240914 385398
rect 244794 710598 245414 711590
rect 244794 710362 244826 710598
rect 245062 710362 245146 710598
rect 245382 710362 245414 710598
rect 244794 710278 245414 710362
rect 244794 710042 244826 710278
rect 245062 710042 245146 710278
rect 245382 710042 245414 710278
rect 244794 678454 245414 710042
rect 244794 678218 244826 678454
rect 245062 678218 245146 678454
rect 245382 678218 245414 678454
rect 244794 678134 245414 678218
rect 244794 677898 244826 678134
rect 245062 677898 245146 678134
rect 245382 677898 245414 678134
rect 244794 642454 245414 677898
rect 244794 642218 244826 642454
rect 245062 642218 245146 642454
rect 245382 642218 245414 642454
rect 244794 642134 245414 642218
rect 244794 641898 244826 642134
rect 245062 641898 245146 642134
rect 245382 641898 245414 642134
rect 244794 606454 245414 641898
rect 244794 606218 244826 606454
rect 245062 606218 245146 606454
rect 245382 606218 245414 606454
rect 244794 606134 245414 606218
rect 244794 605898 244826 606134
rect 245062 605898 245146 606134
rect 245382 605898 245414 606134
rect 244794 570454 245414 605898
rect 244794 570218 244826 570454
rect 245062 570218 245146 570454
rect 245382 570218 245414 570454
rect 244794 570134 245414 570218
rect 244794 569898 244826 570134
rect 245062 569898 245146 570134
rect 245382 569898 245414 570134
rect 244794 534454 245414 569898
rect 244794 534218 244826 534454
rect 245062 534218 245146 534454
rect 245382 534218 245414 534454
rect 244794 534134 245414 534218
rect 244794 533898 244826 534134
rect 245062 533898 245146 534134
rect 245382 533898 245414 534134
rect 244794 498454 245414 533898
rect 244794 498218 244826 498454
rect 245062 498218 245146 498454
rect 245382 498218 245414 498454
rect 244794 498134 245414 498218
rect 244794 497898 244826 498134
rect 245062 497898 245146 498134
rect 245382 497898 245414 498134
rect 244794 462454 245414 497898
rect 244794 462218 244826 462454
rect 245062 462218 245146 462454
rect 245382 462218 245414 462454
rect 244794 462134 245414 462218
rect 244794 461898 244826 462134
rect 245062 461898 245146 462134
rect 245382 461898 245414 462134
rect 244794 426454 245414 461898
rect 244794 426218 244826 426454
rect 245062 426218 245146 426454
rect 245382 426218 245414 426454
rect 244794 426134 245414 426218
rect 244794 425898 244826 426134
rect 245062 425898 245146 426134
rect 245382 425898 245414 426134
rect 244794 390454 245414 425898
rect 244794 390218 244826 390454
rect 245062 390218 245146 390454
rect 245382 390218 245414 390454
rect 244794 390134 245414 390218
rect 244794 389898 244826 390134
rect 245062 389898 245146 390134
rect 245382 389898 245414 390134
rect 244794 384000 245414 389898
rect 249294 711558 249914 711590
rect 249294 711322 249326 711558
rect 249562 711322 249646 711558
rect 249882 711322 249914 711558
rect 249294 711238 249914 711322
rect 249294 711002 249326 711238
rect 249562 711002 249646 711238
rect 249882 711002 249914 711238
rect 249294 682954 249914 711002
rect 249294 682718 249326 682954
rect 249562 682718 249646 682954
rect 249882 682718 249914 682954
rect 249294 682634 249914 682718
rect 249294 682398 249326 682634
rect 249562 682398 249646 682634
rect 249882 682398 249914 682634
rect 249294 646954 249914 682398
rect 249294 646718 249326 646954
rect 249562 646718 249646 646954
rect 249882 646718 249914 646954
rect 249294 646634 249914 646718
rect 249294 646398 249326 646634
rect 249562 646398 249646 646634
rect 249882 646398 249914 646634
rect 249294 610954 249914 646398
rect 249294 610718 249326 610954
rect 249562 610718 249646 610954
rect 249882 610718 249914 610954
rect 249294 610634 249914 610718
rect 249294 610398 249326 610634
rect 249562 610398 249646 610634
rect 249882 610398 249914 610634
rect 249294 574954 249914 610398
rect 249294 574718 249326 574954
rect 249562 574718 249646 574954
rect 249882 574718 249914 574954
rect 249294 574634 249914 574718
rect 249294 574398 249326 574634
rect 249562 574398 249646 574634
rect 249882 574398 249914 574634
rect 249294 538954 249914 574398
rect 249294 538718 249326 538954
rect 249562 538718 249646 538954
rect 249882 538718 249914 538954
rect 249294 538634 249914 538718
rect 249294 538398 249326 538634
rect 249562 538398 249646 538634
rect 249882 538398 249914 538634
rect 249294 502954 249914 538398
rect 249294 502718 249326 502954
rect 249562 502718 249646 502954
rect 249882 502718 249914 502954
rect 249294 502634 249914 502718
rect 249294 502398 249326 502634
rect 249562 502398 249646 502634
rect 249882 502398 249914 502634
rect 249294 466954 249914 502398
rect 249294 466718 249326 466954
rect 249562 466718 249646 466954
rect 249882 466718 249914 466954
rect 249294 466634 249914 466718
rect 249294 466398 249326 466634
rect 249562 466398 249646 466634
rect 249882 466398 249914 466634
rect 249294 430954 249914 466398
rect 249294 430718 249326 430954
rect 249562 430718 249646 430954
rect 249882 430718 249914 430954
rect 249294 430634 249914 430718
rect 249294 430398 249326 430634
rect 249562 430398 249646 430634
rect 249882 430398 249914 430634
rect 249294 394954 249914 430398
rect 249294 394718 249326 394954
rect 249562 394718 249646 394954
rect 249882 394718 249914 394954
rect 249294 394634 249914 394718
rect 249294 394398 249326 394634
rect 249562 394398 249646 394634
rect 249882 394398 249914 394634
rect 249294 384000 249914 394398
rect 253794 704838 254414 711590
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 687454 254414 704282
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 651454 254414 686898
rect 253794 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 254414 651454
rect 253794 651134 254414 651218
rect 253794 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 254414 651134
rect 253794 615454 254414 650898
rect 253794 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 254414 615454
rect 253794 615134 254414 615218
rect 253794 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 254414 615134
rect 253794 579454 254414 614898
rect 253794 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 254414 579454
rect 253794 579134 254414 579218
rect 253794 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 254414 579134
rect 253794 543454 254414 578898
rect 253794 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 254414 543454
rect 253794 543134 254414 543218
rect 253794 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 254414 543134
rect 253794 507454 254414 542898
rect 253794 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 254414 507454
rect 253794 507134 254414 507218
rect 253794 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 254414 507134
rect 253794 471454 254414 506898
rect 253794 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 254414 471454
rect 253794 471134 254414 471218
rect 253794 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 254414 471134
rect 253794 435454 254414 470898
rect 253794 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 254414 435454
rect 253794 435134 254414 435218
rect 253794 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 254414 435134
rect 253794 399454 254414 434898
rect 253794 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 254414 399454
rect 253794 399134 254414 399218
rect 253794 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 254414 399134
rect 253794 384000 254414 398898
rect 258294 705798 258914 711590
rect 258294 705562 258326 705798
rect 258562 705562 258646 705798
rect 258882 705562 258914 705798
rect 258294 705478 258914 705562
rect 258294 705242 258326 705478
rect 258562 705242 258646 705478
rect 258882 705242 258914 705478
rect 258294 691954 258914 705242
rect 258294 691718 258326 691954
rect 258562 691718 258646 691954
rect 258882 691718 258914 691954
rect 258294 691634 258914 691718
rect 258294 691398 258326 691634
rect 258562 691398 258646 691634
rect 258882 691398 258914 691634
rect 258294 655954 258914 691398
rect 258294 655718 258326 655954
rect 258562 655718 258646 655954
rect 258882 655718 258914 655954
rect 258294 655634 258914 655718
rect 258294 655398 258326 655634
rect 258562 655398 258646 655634
rect 258882 655398 258914 655634
rect 258294 619954 258914 655398
rect 258294 619718 258326 619954
rect 258562 619718 258646 619954
rect 258882 619718 258914 619954
rect 258294 619634 258914 619718
rect 258294 619398 258326 619634
rect 258562 619398 258646 619634
rect 258882 619398 258914 619634
rect 258294 583954 258914 619398
rect 258294 583718 258326 583954
rect 258562 583718 258646 583954
rect 258882 583718 258914 583954
rect 258294 583634 258914 583718
rect 258294 583398 258326 583634
rect 258562 583398 258646 583634
rect 258882 583398 258914 583634
rect 258294 547954 258914 583398
rect 258294 547718 258326 547954
rect 258562 547718 258646 547954
rect 258882 547718 258914 547954
rect 258294 547634 258914 547718
rect 258294 547398 258326 547634
rect 258562 547398 258646 547634
rect 258882 547398 258914 547634
rect 258294 511954 258914 547398
rect 258294 511718 258326 511954
rect 258562 511718 258646 511954
rect 258882 511718 258914 511954
rect 258294 511634 258914 511718
rect 258294 511398 258326 511634
rect 258562 511398 258646 511634
rect 258882 511398 258914 511634
rect 258294 475954 258914 511398
rect 258294 475718 258326 475954
rect 258562 475718 258646 475954
rect 258882 475718 258914 475954
rect 258294 475634 258914 475718
rect 258294 475398 258326 475634
rect 258562 475398 258646 475634
rect 258882 475398 258914 475634
rect 258294 439954 258914 475398
rect 258294 439718 258326 439954
rect 258562 439718 258646 439954
rect 258882 439718 258914 439954
rect 258294 439634 258914 439718
rect 258294 439398 258326 439634
rect 258562 439398 258646 439634
rect 258882 439398 258914 439634
rect 258294 403954 258914 439398
rect 258294 403718 258326 403954
rect 258562 403718 258646 403954
rect 258882 403718 258914 403954
rect 258294 403634 258914 403718
rect 258294 403398 258326 403634
rect 258562 403398 258646 403634
rect 258882 403398 258914 403634
rect 258294 384000 258914 403398
rect 262794 706758 263414 711590
rect 262794 706522 262826 706758
rect 263062 706522 263146 706758
rect 263382 706522 263414 706758
rect 262794 706438 263414 706522
rect 262794 706202 262826 706438
rect 263062 706202 263146 706438
rect 263382 706202 263414 706438
rect 262794 696454 263414 706202
rect 262794 696218 262826 696454
rect 263062 696218 263146 696454
rect 263382 696218 263414 696454
rect 262794 696134 263414 696218
rect 262794 695898 262826 696134
rect 263062 695898 263146 696134
rect 263382 695898 263414 696134
rect 262794 660454 263414 695898
rect 262794 660218 262826 660454
rect 263062 660218 263146 660454
rect 263382 660218 263414 660454
rect 262794 660134 263414 660218
rect 262794 659898 262826 660134
rect 263062 659898 263146 660134
rect 263382 659898 263414 660134
rect 262794 624454 263414 659898
rect 262794 624218 262826 624454
rect 263062 624218 263146 624454
rect 263382 624218 263414 624454
rect 262794 624134 263414 624218
rect 262794 623898 262826 624134
rect 263062 623898 263146 624134
rect 263382 623898 263414 624134
rect 262794 588454 263414 623898
rect 262794 588218 262826 588454
rect 263062 588218 263146 588454
rect 263382 588218 263414 588454
rect 262794 588134 263414 588218
rect 262794 587898 262826 588134
rect 263062 587898 263146 588134
rect 263382 587898 263414 588134
rect 262794 552454 263414 587898
rect 262794 552218 262826 552454
rect 263062 552218 263146 552454
rect 263382 552218 263414 552454
rect 262794 552134 263414 552218
rect 262794 551898 262826 552134
rect 263062 551898 263146 552134
rect 263382 551898 263414 552134
rect 262794 516454 263414 551898
rect 262794 516218 262826 516454
rect 263062 516218 263146 516454
rect 263382 516218 263414 516454
rect 262794 516134 263414 516218
rect 262794 515898 262826 516134
rect 263062 515898 263146 516134
rect 263382 515898 263414 516134
rect 262794 480454 263414 515898
rect 262794 480218 262826 480454
rect 263062 480218 263146 480454
rect 263382 480218 263414 480454
rect 262794 480134 263414 480218
rect 262794 479898 262826 480134
rect 263062 479898 263146 480134
rect 263382 479898 263414 480134
rect 262794 444454 263414 479898
rect 262794 444218 262826 444454
rect 263062 444218 263146 444454
rect 263382 444218 263414 444454
rect 262794 444134 263414 444218
rect 262794 443898 262826 444134
rect 263062 443898 263146 444134
rect 263382 443898 263414 444134
rect 262794 408454 263414 443898
rect 262794 408218 262826 408454
rect 263062 408218 263146 408454
rect 263382 408218 263414 408454
rect 262794 408134 263414 408218
rect 262794 407898 262826 408134
rect 263062 407898 263146 408134
rect 263382 407898 263414 408134
rect 262794 384000 263414 407898
rect 267294 707718 267914 711590
rect 267294 707482 267326 707718
rect 267562 707482 267646 707718
rect 267882 707482 267914 707718
rect 267294 707398 267914 707482
rect 267294 707162 267326 707398
rect 267562 707162 267646 707398
rect 267882 707162 267914 707398
rect 267294 700954 267914 707162
rect 267294 700718 267326 700954
rect 267562 700718 267646 700954
rect 267882 700718 267914 700954
rect 267294 700634 267914 700718
rect 267294 700398 267326 700634
rect 267562 700398 267646 700634
rect 267882 700398 267914 700634
rect 267294 664954 267914 700398
rect 267294 664718 267326 664954
rect 267562 664718 267646 664954
rect 267882 664718 267914 664954
rect 267294 664634 267914 664718
rect 267294 664398 267326 664634
rect 267562 664398 267646 664634
rect 267882 664398 267914 664634
rect 267294 628954 267914 664398
rect 267294 628718 267326 628954
rect 267562 628718 267646 628954
rect 267882 628718 267914 628954
rect 267294 628634 267914 628718
rect 267294 628398 267326 628634
rect 267562 628398 267646 628634
rect 267882 628398 267914 628634
rect 267294 592954 267914 628398
rect 267294 592718 267326 592954
rect 267562 592718 267646 592954
rect 267882 592718 267914 592954
rect 267294 592634 267914 592718
rect 267294 592398 267326 592634
rect 267562 592398 267646 592634
rect 267882 592398 267914 592634
rect 267294 556954 267914 592398
rect 267294 556718 267326 556954
rect 267562 556718 267646 556954
rect 267882 556718 267914 556954
rect 267294 556634 267914 556718
rect 267294 556398 267326 556634
rect 267562 556398 267646 556634
rect 267882 556398 267914 556634
rect 267294 520954 267914 556398
rect 267294 520718 267326 520954
rect 267562 520718 267646 520954
rect 267882 520718 267914 520954
rect 267294 520634 267914 520718
rect 267294 520398 267326 520634
rect 267562 520398 267646 520634
rect 267882 520398 267914 520634
rect 267294 484954 267914 520398
rect 267294 484718 267326 484954
rect 267562 484718 267646 484954
rect 267882 484718 267914 484954
rect 267294 484634 267914 484718
rect 267294 484398 267326 484634
rect 267562 484398 267646 484634
rect 267882 484398 267914 484634
rect 267294 448954 267914 484398
rect 267294 448718 267326 448954
rect 267562 448718 267646 448954
rect 267882 448718 267914 448954
rect 267294 448634 267914 448718
rect 267294 448398 267326 448634
rect 267562 448398 267646 448634
rect 267882 448398 267914 448634
rect 267294 412954 267914 448398
rect 267294 412718 267326 412954
rect 267562 412718 267646 412954
rect 267882 412718 267914 412954
rect 267294 412634 267914 412718
rect 267294 412398 267326 412634
rect 267562 412398 267646 412634
rect 267882 412398 267914 412634
rect 267294 384000 267914 412398
rect 271794 708678 272414 711590
rect 271794 708442 271826 708678
rect 272062 708442 272146 708678
rect 272382 708442 272414 708678
rect 271794 708358 272414 708442
rect 271794 708122 271826 708358
rect 272062 708122 272146 708358
rect 272382 708122 272414 708358
rect 271794 669454 272414 708122
rect 271794 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 272414 669454
rect 271794 669134 272414 669218
rect 271794 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 272414 669134
rect 271794 633454 272414 668898
rect 271794 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 272414 633454
rect 271794 633134 272414 633218
rect 271794 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 272414 633134
rect 271794 597454 272414 632898
rect 271794 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 272414 597454
rect 271794 597134 272414 597218
rect 271794 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 272414 597134
rect 271794 561454 272414 596898
rect 271794 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 272414 561454
rect 271794 561134 272414 561218
rect 271794 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 272414 561134
rect 271794 525454 272414 560898
rect 271794 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 272414 525454
rect 271794 525134 272414 525218
rect 271794 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 272414 525134
rect 271794 489454 272414 524898
rect 271794 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 272414 489454
rect 271794 489134 272414 489218
rect 271794 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 272414 489134
rect 271794 453454 272414 488898
rect 271794 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 272414 453454
rect 271794 453134 272414 453218
rect 271794 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 272414 453134
rect 271794 417454 272414 452898
rect 271794 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 272414 417454
rect 271794 417134 272414 417218
rect 271794 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 272414 417134
rect 271794 384000 272414 416898
rect 276294 709638 276914 711590
rect 276294 709402 276326 709638
rect 276562 709402 276646 709638
rect 276882 709402 276914 709638
rect 276294 709318 276914 709402
rect 276294 709082 276326 709318
rect 276562 709082 276646 709318
rect 276882 709082 276914 709318
rect 276294 673954 276914 709082
rect 276294 673718 276326 673954
rect 276562 673718 276646 673954
rect 276882 673718 276914 673954
rect 276294 673634 276914 673718
rect 276294 673398 276326 673634
rect 276562 673398 276646 673634
rect 276882 673398 276914 673634
rect 276294 637954 276914 673398
rect 276294 637718 276326 637954
rect 276562 637718 276646 637954
rect 276882 637718 276914 637954
rect 276294 637634 276914 637718
rect 276294 637398 276326 637634
rect 276562 637398 276646 637634
rect 276882 637398 276914 637634
rect 276294 601954 276914 637398
rect 276294 601718 276326 601954
rect 276562 601718 276646 601954
rect 276882 601718 276914 601954
rect 276294 601634 276914 601718
rect 276294 601398 276326 601634
rect 276562 601398 276646 601634
rect 276882 601398 276914 601634
rect 276294 565954 276914 601398
rect 276294 565718 276326 565954
rect 276562 565718 276646 565954
rect 276882 565718 276914 565954
rect 276294 565634 276914 565718
rect 276294 565398 276326 565634
rect 276562 565398 276646 565634
rect 276882 565398 276914 565634
rect 276294 529954 276914 565398
rect 276294 529718 276326 529954
rect 276562 529718 276646 529954
rect 276882 529718 276914 529954
rect 276294 529634 276914 529718
rect 276294 529398 276326 529634
rect 276562 529398 276646 529634
rect 276882 529398 276914 529634
rect 276294 493954 276914 529398
rect 276294 493718 276326 493954
rect 276562 493718 276646 493954
rect 276882 493718 276914 493954
rect 276294 493634 276914 493718
rect 276294 493398 276326 493634
rect 276562 493398 276646 493634
rect 276882 493398 276914 493634
rect 276294 457954 276914 493398
rect 276294 457718 276326 457954
rect 276562 457718 276646 457954
rect 276882 457718 276914 457954
rect 276294 457634 276914 457718
rect 276294 457398 276326 457634
rect 276562 457398 276646 457634
rect 276882 457398 276914 457634
rect 276294 421954 276914 457398
rect 276294 421718 276326 421954
rect 276562 421718 276646 421954
rect 276882 421718 276914 421954
rect 276294 421634 276914 421718
rect 276294 421398 276326 421634
rect 276562 421398 276646 421634
rect 276882 421398 276914 421634
rect 276294 385954 276914 421398
rect 276294 385718 276326 385954
rect 276562 385718 276646 385954
rect 276882 385718 276914 385954
rect 276294 385634 276914 385718
rect 276294 385398 276326 385634
rect 276562 385398 276646 385634
rect 276882 385398 276914 385634
rect 276294 384000 276914 385398
rect 280794 710598 281414 711590
rect 280794 710362 280826 710598
rect 281062 710362 281146 710598
rect 281382 710362 281414 710598
rect 280794 710278 281414 710362
rect 280794 710042 280826 710278
rect 281062 710042 281146 710278
rect 281382 710042 281414 710278
rect 280794 678454 281414 710042
rect 280794 678218 280826 678454
rect 281062 678218 281146 678454
rect 281382 678218 281414 678454
rect 280794 678134 281414 678218
rect 280794 677898 280826 678134
rect 281062 677898 281146 678134
rect 281382 677898 281414 678134
rect 280794 642454 281414 677898
rect 280794 642218 280826 642454
rect 281062 642218 281146 642454
rect 281382 642218 281414 642454
rect 280794 642134 281414 642218
rect 280794 641898 280826 642134
rect 281062 641898 281146 642134
rect 281382 641898 281414 642134
rect 280794 606454 281414 641898
rect 280794 606218 280826 606454
rect 281062 606218 281146 606454
rect 281382 606218 281414 606454
rect 280794 606134 281414 606218
rect 280794 605898 280826 606134
rect 281062 605898 281146 606134
rect 281382 605898 281414 606134
rect 280794 570454 281414 605898
rect 280794 570218 280826 570454
rect 281062 570218 281146 570454
rect 281382 570218 281414 570454
rect 280794 570134 281414 570218
rect 280794 569898 280826 570134
rect 281062 569898 281146 570134
rect 281382 569898 281414 570134
rect 280794 534454 281414 569898
rect 280794 534218 280826 534454
rect 281062 534218 281146 534454
rect 281382 534218 281414 534454
rect 280794 534134 281414 534218
rect 280794 533898 280826 534134
rect 281062 533898 281146 534134
rect 281382 533898 281414 534134
rect 280794 498454 281414 533898
rect 280794 498218 280826 498454
rect 281062 498218 281146 498454
rect 281382 498218 281414 498454
rect 280794 498134 281414 498218
rect 280794 497898 280826 498134
rect 281062 497898 281146 498134
rect 281382 497898 281414 498134
rect 280794 462454 281414 497898
rect 280794 462218 280826 462454
rect 281062 462218 281146 462454
rect 281382 462218 281414 462454
rect 280794 462134 281414 462218
rect 280794 461898 280826 462134
rect 281062 461898 281146 462134
rect 281382 461898 281414 462134
rect 280794 426454 281414 461898
rect 280794 426218 280826 426454
rect 281062 426218 281146 426454
rect 281382 426218 281414 426454
rect 280794 426134 281414 426218
rect 280794 425898 280826 426134
rect 281062 425898 281146 426134
rect 281382 425898 281414 426134
rect 280794 390454 281414 425898
rect 280794 390218 280826 390454
rect 281062 390218 281146 390454
rect 281382 390218 281414 390454
rect 280794 390134 281414 390218
rect 280794 389898 280826 390134
rect 281062 389898 281146 390134
rect 281382 389898 281414 390134
rect 280794 384000 281414 389898
rect 285294 711558 285914 711590
rect 285294 711322 285326 711558
rect 285562 711322 285646 711558
rect 285882 711322 285914 711558
rect 285294 711238 285914 711322
rect 285294 711002 285326 711238
rect 285562 711002 285646 711238
rect 285882 711002 285914 711238
rect 285294 682954 285914 711002
rect 285294 682718 285326 682954
rect 285562 682718 285646 682954
rect 285882 682718 285914 682954
rect 285294 682634 285914 682718
rect 285294 682398 285326 682634
rect 285562 682398 285646 682634
rect 285882 682398 285914 682634
rect 285294 646954 285914 682398
rect 285294 646718 285326 646954
rect 285562 646718 285646 646954
rect 285882 646718 285914 646954
rect 285294 646634 285914 646718
rect 285294 646398 285326 646634
rect 285562 646398 285646 646634
rect 285882 646398 285914 646634
rect 285294 610954 285914 646398
rect 285294 610718 285326 610954
rect 285562 610718 285646 610954
rect 285882 610718 285914 610954
rect 285294 610634 285914 610718
rect 285294 610398 285326 610634
rect 285562 610398 285646 610634
rect 285882 610398 285914 610634
rect 285294 574954 285914 610398
rect 285294 574718 285326 574954
rect 285562 574718 285646 574954
rect 285882 574718 285914 574954
rect 285294 574634 285914 574718
rect 285294 574398 285326 574634
rect 285562 574398 285646 574634
rect 285882 574398 285914 574634
rect 285294 538954 285914 574398
rect 285294 538718 285326 538954
rect 285562 538718 285646 538954
rect 285882 538718 285914 538954
rect 285294 538634 285914 538718
rect 285294 538398 285326 538634
rect 285562 538398 285646 538634
rect 285882 538398 285914 538634
rect 285294 502954 285914 538398
rect 285294 502718 285326 502954
rect 285562 502718 285646 502954
rect 285882 502718 285914 502954
rect 285294 502634 285914 502718
rect 285294 502398 285326 502634
rect 285562 502398 285646 502634
rect 285882 502398 285914 502634
rect 285294 466954 285914 502398
rect 285294 466718 285326 466954
rect 285562 466718 285646 466954
rect 285882 466718 285914 466954
rect 285294 466634 285914 466718
rect 285294 466398 285326 466634
rect 285562 466398 285646 466634
rect 285882 466398 285914 466634
rect 285294 430954 285914 466398
rect 285294 430718 285326 430954
rect 285562 430718 285646 430954
rect 285882 430718 285914 430954
rect 285294 430634 285914 430718
rect 285294 430398 285326 430634
rect 285562 430398 285646 430634
rect 285882 430398 285914 430634
rect 285294 394954 285914 430398
rect 285294 394718 285326 394954
rect 285562 394718 285646 394954
rect 285882 394718 285914 394954
rect 285294 394634 285914 394718
rect 285294 394398 285326 394634
rect 285562 394398 285646 394634
rect 285882 394398 285914 394634
rect 285294 384000 285914 394398
rect 289794 704838 290414 711590
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 651454 290414 686898
rect 289794 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 290414 651454
rect 289794 651134 290414 651218
rect 289794 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 290414 651134
rect 289794 615454 290414 650898
rect 289794 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 290414 615454
rect 289794 615134 290414 615218
rect 289794 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 290414 615134
rect 289794 579454 290414 614898
rect 289794 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 290414 579454
rect 289794 579134 290414 579218
rect 289794 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 290414 579134
rect 289794 543454 290414 578898
rect 289794 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 290414 543454
rect 289794 543134 290414 543218
rect 289794 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 290414 543134
rect 289794 507454 290414 542898
rect 289794 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 290414 507454
rect 289794 507134 290414 507218
rect 289794 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 290414 507134
rect 289794 471454 290414 506898
rect 289794 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 290414 471454
rect 289794 471134 290414 471218
rect 289794 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 290414 471134
rect 289794 435454 290414 470898
rect 289794 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 290414 435454
rect 289794 435134 290414 435218
rect 289794 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 290414 435134
rect 289794 399454 290414 434898
rect 289794 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 290414 399454
rect 289794 399134 290414 399218
rect 289794 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 290414 399134
rect 289794 384000 290414 398898
rect 294294 705798 294914 711590
rect 294294 705562 294326 705798
rect 294562 705562 294646 705798
rect 294882 705562 294914 705798
rect 294294 705478 294914 705562
rect 294294 705242 294326 705478
rect 294562 705242 294646 705478
rect 294882 705242 294914 705478
rect 294294 691954 294914 705242
rect 294294 691718 294326 691954
rect 294562 691718 294646 691954
rect 294882 691718 294914 691954
rect 294294 691634 294914 691718
rect 294294 691398 294326 691634
rect 294562 691398 294646 691634
rect 294882 691398 294914 691634
rect 294294 655954 294914 691398
rect 294294 655718 294326 655954
rect 294562 655718 294646 655954
rect 294882 655718 294914 655954
rect 294294 655634 294914 655718
rect 294294 655398 294326 655634
rect 294562 655398 294646 655634
rect 294882 655398 294914 655634
rect 294294 619954 294914 655398
rect 294294 619718 294326 619954
rect 294562 619718 294646 619954
rect 294882 619718 294914 619954
rect 294294 619634 294914 619718
rect 294294 619398 294326 619634
rect 294562 619398 294646 619634
rect 294882 619398 294914 619634
rect 294294 583954 294914 619398
rect 294294 583718 294326 583954
rect 294562 583718 294646 583954
rect 294882 583718 294914 583954
rect 294294 583634 294914 583718
rect 294294 583398 294326 583634
rect 294562 583398 294646 583634
rect 294882 583398 294914 583634
rect 294294 547954 294914 583398
rect 294294 547718 294326 547954
rect 294562 547718 294646 547954
rect 294882 547718 294914 547954
rect 294294 547634 294914 547718
rect 294294 547398 294326 547634
rect 294562 547398 294646 547634
rect 294882 547398 294914 547634
rect 294294 511954 294914 547398
rect 294294 511718 294326 511954
rect 294562 511718 294646 511954
rect 294882 511718 294914 511954
rect 294294 511634 294914 511718
rect 294294 511398 294326 511634
rect 294562 511398 294646 511634
rect 294882 511398 294914 511634
rect 294294 475954 294914 511398
rect 294294 475718 294326 475954
rect 294562 475718 294646 475954
rect 294882 475718 294914 475954
rect 294294 475634 294914 475718
rect 294294 475398 294326 475634
rect 294562 475398 294646 475634
rect 294882 475398 294914 475634
rect 294294 439954 294914 475398
rect 294294 439718 294326 439954
rect 294562 439718 294646 439954
rect 294882 439718 294914 439954
rect 294294 439634 294914 439718
rect 294294 439398 294326 439634
rect 294562 439398 294646 439634
rect 294882 439398 294914 439634
rect 294294 403954 294914 439398
rect 294294 403718 294326 403954
rect 294562 403718 294646 403954
rect 294882 403718 294914 403954
rect 294294 403634 294914 403718
rect 294294 403398 294326 403634
rect 294562 403398 294646 403634
rect 294882 403398 294914 403634
rect 293355 384844 293421 384845
rect 293355 384780 293356 384844
rect 293420 384780 293421 384844
rect 293355 384779 293421 384780
rect 290779 384436 290845 384437
rect 290779 384372 290780 384436
rect 290844 384372 290845 384436
rect 290779 384371 290845 384372
rect 290595 382940 290661 382941
rect 290595 382876 290596 382940
rect 290660 382876 290661 382940
rect 290595 382875 290661 382876
rect 283971 382124 284037 382125
rect 283971 382060 283972 382124
rect 284036 382060 284037 382124
rect 283971 382059 284037 382060
rect 258763 381852 258829 381853
rect 258763 381788 258764 381852
rect 258828 381788 258829 381852
rect 258763 381787 258829 381788
rect 273851 381852 273917 381853
rect 273851 381788 273852 381852
rect 273916 381788 273917 381852
rect 273851 381787 273917 381788
rect 276059 381852 276125 381853
rect 276059 381788 276060 381852
rect 276124 381788 276125 381852
rect 276059 381787 276125 381788
rect 280291 381852 280357 381853
rect 280291 381788 280292 381852
rect 280356 381788 280357 381852
rect 280291 381787 280357 381788
rect 282499 381852 282565 381853
rect 282499 381788 282500 381852
rect 282564 381788 282565 381852
rect 282499 381787 282565 381788
rect 239995 381444 240061 381445
rect 239995 381380 239996 381444
rect 240060 381380 240061 381444
rect 239995 381379 240061 381380
rect 242387 381444 242453 381445
rect 242387 381380 242388 381444
rect 242452 381380 242453 381444
rect 242387 381379 242453 381380
rect 245515 381444 245581 381445
rect 245515 381380 245516 381444
rect 245580 381380 245581 381444
rect 245515 381379 245581 381380
rect 239998 380221 240058 381379
rect 242390 381037 242450 381379
rect 242387 381036 242453 381037
rect 242387 380972 242388 381036
rect 242452 380972 242453 381036
rect 242387 380971 242453 380972
rect 245518 380357 245578 381379
rect 258766 381173 258826 381787
rect 258763 381172 258829 381173
rect 258763 381108 258764 381172
rect 258828 381108 258829 381172
rect 258763 381107 258829 381108
rect 273854 380629 273914 381787
rect 273851 380628 273917 380629
rect 273851 380564 273852 380628
rect 273916 380564 273917 380628
rect 273851 380563 273917 380564
rect 276062 380493 276122 381787
rect 280294 381173 280354 381787
rect 280291 381172 280357 381173
rect 280291 381108 280292 381172
rect 280356 381108 280357 381172
rect 280291 381107 280357 381108
rect 282502 380493 282562 381787
rect 283974 380629 284034 382059
rect 288755 381988 288821 381989
rect 288755 381924 288756 381988
rect 288820 381924 288821 381988
rect 288755 381923 288821 381924
rect 288939 381988 289005 381989
rect 288939 381924 288940 381988
rect 289004 381924 289005 381988
rect 288939 381923 289005 381924
rect 283971 380628 284037 380629
rect 283971 380564 283972 380628
rect 284036 380564 284037 380628
rect 283971 380563 284037 380564
rect 276059 380492 276125 380493
rect 276059 380428 276060 380492
rect 276124 380428 276125 380492
rect 276059 380427 276125 380428
rect 282499 380492 282565 380493
rect 282499 380428 282500 380492
rect 282564 380428 282565 380492
rect 282499 380427 282565 380428
rect 245515 380356 245581 380357
rect 245515 380292 245516 380356
rect 245580 380292 245581 380356
rect 245515 380291 245581 380292
rect 239995 380220 240061 380221
rect 239995 380156 239996 380220
rect 240060 380156 240061 380220
rect 239995 380155 240061 380156
rect 254568 367954 254888 367986
rect 254568 367718 254610 367954
rect 254846 367718 254888 367954
rect 254568 367634 254888 367718
rect 254568 367398 254610 367634
rect 254846 367398 254888 367634
rect 254568 367366 254888 367398
rect 285288 367954 285608 367986
rect 285288 367718 285330 367954
rect 285566 367718 285608 367954
rect 285288 367634 285608 367718
rect 285288 367398 285330 367634
rect 285566 367398 285608 367634
rect 285288 367366 285608 367398
rect 269928 363454 270248 363486
rect 269928 363218 269970 363454
rect 270206 363218 270248 363454
rect 269928 363134 270248 363218
rect 269928 362898 269970 363134
rect 270206 362898 270248 363134
rect 269928 362866 270248 362898
rect 238891 339964 238957 339965
rect 238891 339900 238892 339964
rect 238956 339900 238957 339964
rect 238891 339899 238957 339900
rect 239627 339964 239693 339965
rect 239627 339900 239628 339964
rect 239692 339900 239693 339964
rect 239627 339899 239693 339900
rect 245883 338196 245949 338197
rect 245883 338132 245884 338196
rect 245948 338132 245949 338196
rect 245883 338131 245949 338132
rect 254531 338196 254597 338197
rect 254531 338132 254532 338196
rect 254596 338132 254597 338196
rect 254531 338131 254597 338132
rect 255635 338196 255701 338197
rect 255635 338132 255636 338196
rect 255700 338132 255701 338196
rect 255635 338131 255701 338132
rect 245699 337924 245765 337925
rect 245699 337860 245700 337924
rect 245764 337860 245765 337924
rect 245699 337859 245765 337860
rect 240294 313954 240914 336000
rect 243491 335340 243557 335341
rect 243491 335276 243492 335340
rect 243556 335276 243557 335340
rect 243491 335275 243557 335276
rect 240294 313718 240326 313954
rect 240562 313718 240646 313954
rect 240882 313718 240914 313954
rect 240294 313634 240914 313718
rect 240294 313398 240326 313634
rect 240562 313398 240646 313634
rect 240882 313398 240914 313634
rect 240294 277954 240914 313398
rect 240294 277718 240326 277954
rect 240562 277718 240646 277954
rect 240882 277718 240914 277954
rect 240294 277634 240914 277718
rect 240294 277398 240326 277634
rect 240562 277398 240646 277634
rect 240882 277398 240914 277634
rect 240294 241954 240914 277398
rect 240294 241718 240326 241954
rect 240562 241718 240646 241954
rect 240882 241718 240914 241954
rect 240294 241634 240914 241718
rect 240294 241398 240326 241634
rect 240562 241398 240646 241634
rect 240882 241398 240914 241634
rect 240294 205954 240914 241398
rect 240294 205718 240326 205954
rect 240562 205718 240646 205954
rect 240882 205718 240914 205954
rect 240294 205634 240914 205718
rect 240294 205398 240326 205634
rect 240562 205398 240646 205634
rect 240882 205398 240914 205634
rect 240294 169954 240914 205398
rect 240294 169718 240326 169954
rect 240562 169718 240646 169954
rect 240882 169718 240914 169954
rect 240294 169634 240914 169718
rect 240294 169398 240326 169634
rect 240562 169398 240646 169634
rect 240882 169398 240914 169634
rect 240294 133954 240914 169398
rect 240294 133718 240326 133954
rect 240562 133718 240646 133954
rect 240882 133718 240914 133954
rect 240294 133634 240914 133718
rect 240294 133398 240326 133634
rect 240562 133398 240646 133634
rect 240882 133398 240914 133634
rect 238523 107676 238589 107677
rect 238523 107612 238524 107676
rect 238588 107612 238589 107676
rect 238523 107611 238589 107612
rect 240294 97954 240914 133398
rect 238339 97748 238405 97749
rect 238339 97684 238340 97748
rect 238404 97684 238405 97748
rect 238339 97683 238405 97684
rect 240294 97718 240326 97954
rect 240562 97718 240646 97954
rect 240882 97718 240914 97954
rect 240294 97634 240914 97718
rect 237235 97612 237301 97613
rect 237235 97548 237236 97612
rect 237300 97548 237301 97612
rect 237235 97547 237301 97548
rect 235794 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 236414 93454
rect 235794 93134 236414 93218
rect 235794 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 236414 93134
rect 235794 57454 236414 92898
rect 235794 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 236414 57454
rect 235794 57134 236414 57218
rect 235794 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 236414 57134
rect 235794 21454 236414 56898
rect 235794 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 236414 21454
rect 235794 21134 236414 21218
rect 235794 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 236414 21134
rect 235794 -4186 236414 20898
rect 235794 -4422 235826 -4186
rect 236062 -4422 236146 -4186
rect 236382 -4422 236414 -4186
rect 235794 -4506 236414 -4422
rect 235794 -4742 235826 -4506
rect 236062 -4742 236146 -4506
rect 236382 -4742 236414 -4506
rect 235794 -7654 236414 -4742
rect 240294 97398 240326 97634
rect 240562 97398 240646 97634
rect 240882 97398 240914 97634
rect 240294 61954 240914 97398
rect 240294 61718 240326 61954
rect 240562 61718 240646 61954
rect 240882 61718 240914 61954
rect 240294 61634 240914 61718
rect 240294 61398 240326 61634
rect 240562 61398 240646 61634
rect 240882 61398 240914 61634
rect 240294 25954 240914 61398
rect 240294 25718 240326 25954
rect 240562 25718 240646 25954
rect 240882 25718 240914 25954
rect 240294 25634 240914 25718
rect 240294 25398 240326 25634
rect 240562 25398 240646 25634
rect 240882 25398 240914 25634
rect 240294 -5146 240914 25398
rect 243494 3365 243554 335275
rect 244794 318454 245414 336000
rect 244794 318218 244826 318454
rect 245062 318218 245146 318454
rect 245382 318218 245414 318454
rect 244794 318134 245414 318218
rect 244794 317898 244826 318134
rect 245062 317898 245146 318134
rect 245382 317898 245414 318134
rect 244794 282454 245414 317898
rect 244794 282218 244826 282454
rect 245062 282218 245146 282454
rect 245382 282218 245414 282454
rect 244794 282134 245414 282218
rect 244794 281898 244826 282134
rect 245062 281898 245146 282134
rect 245382 281898 245414 282134
rect 244794 246454 245414 281898
rect 244794 246218 244826 246454
rect 245062 246218 245146 246454
rect 245382 246218 245414 246454
rect 244794 246134 245414 246218
rect 244794 245898 244826 246134
rect 245062 245898 245146 246134
rect 245382 245898 245414 246134
rect 244794 210454 245414 245898
rect 244794 210218 244826 210454
rect 245062 210218 245146 210454
rect 245382 210218 245414 210454
rect 244794 210134 245414 210218
rect 244794 209898 244826 210134
rect 245062 209898 245146 210134
rect 245382 209898 245414 210134
rect 244794 174454 245414 209898
rect 244794 174218 244826 174454
rect 245062 174218 245146 174454
rect 245382 174218 245414 174454
rect 244794 174134 245414 174218
rect 244794 173898 244826 174134
rect 245062 173898 245146 174134
rect 245382 173898 245414 174134
rect 244794 138454 245414 173898
rect 244794 138218 244826 138454
rect 245062 138218 245146 138454
rect 245382 138218 245414 138454
rect 244794 138134 245414 138218
rect 244794 137898 244826 138134
rect 245062 137898 245146 138134
rect 245382 137898 245414 138134
rect 244794 102454 245414 137898
rect 244794 102218 244826 102454
rect 245062 102218 245146 102454
rect 245382 102218 245414 102454
rect 244794 102134 245414 102218
rect 244794 101898 244826 102134
rect 245062 101898 245146 102134
rect 245382 101898 245414 102134
rect 244794 66454 245414 101898
rect 244794 66218 244826 66454
rect 245062 66218 245146 66454
rect 245382 66218 245414 66454
rect 244794 66134 245414 66218
rect 244794 65898 244826 66134
rect 245062 65898 245146 66134
rect 245382 65898 245414 66134
rect 244794 30454 245414 65898
rect 244794 30218 244826 30454
rect 245062 30218 245146 30454
rect 245382 30218 245414 30454
rect 244794 30134 245414 30218
rect 244794 29898 244826 30134
rect 245062 29898 245146 30134
rect 245382 29898 245414 30134
rect 243491 3364 243557 3365
rect 243491 3300 243492 3364
rect 243556 3300 243557 3364
rect 243491 3299 243557 3300
rect 240294 -5382 240326 -5146
rect 240562 -5382 240646 -5146
rect 240882 -5382 240914 -5146
rect 240294 -5466 240914 -5382
rect 240294 -5702 240326 -5466
rect 240562 -5702 240646 -5466
rect 240882 -5702 240914 -5466
rect 240294 -7654 240914 -5702
rect 244794 -6106 245414 29898
rect 245702 4861 245762 337859
rect 245886 13021 245946 338131
rect 247171 337924 247237 337925
rect 247171 337860 247172 337924
rect 247236 337860 247237 337924
rect 247171 337859 247237 337860
rect 248275 337924 248341 337925
rect 248275 337860 248276 337924
rect 248340 337860 248341 337924
rect 248275 337859 248341 337860
rect 250115 337924 250181 337925
rect 250115 337860 250116 337924
rect 250180 337860 250181 337924
rect 250115 337859 250181 337860
rect 251403 337924 251469 337925
rect 251403 337860 251404 337924
rect 251468 337860 251469 337924
rect 251403 337859 251469 337860
rect 251771 337924 251837 337925
rect 251771 337860 251772 337924
rect 251836 337860 251837 337924
rect 251771 337859 251837 337860
rect 252875 337924 252941 337925
rect 252875 337860 252876 337924
rect 252940 337860 252941 337924
rect 252875 337859 252941 337860
rect 254163 337924 254229 337925
rect 254163 337860 254164 337924
rect 254228 337860 254229 337924
rect 254163 337859 254229 337860
rect 246251 337788 246317 337789
rect 246251 337724 246252 337788
rect 246316 337724 246317 337788
rect 246251 337723 246317 337724
rect 246067 334796 246133 334797
rect 246067 334732 246068 334796
rect 246132 334732 246133 334796
rect 246067 334731 246133 334732
rect 246070 326365 246130 334731
rect 246254 327725 246314 337723
rect 246251 327724 246317 327725
rect 246251 327660 246252 327724
rect 246316 327660 246317 327724
rect 246251 327659 246317 327660
rect 246067 326364 246133 326365
rect 246067 326300 246068 326364
rect 246132 326300 246133 326364
rect 246067 326299 246133 326300
rect 247174 79389 247234 337859
rect 247355 337788 247421 337789
rect 247355 337724 247356 337788
rect 247420 337724 247421 337788
rect 247355 337723 247421 337724
rect 247171 79388 247237 79389
rect 247171 79324 247172 79388
rect 247236 79324 247237 79388
rect 247171 79323 247237 79324
rect 247358 13157 247418 337723
rect 248278 335613 248338 337859
rect 248275 335612 248341 335613
rect 248275 335548 248276 335612
rect 248340 335548 248341 335612
rect 248275 335547 248341 335548
rect 248643 333300 248709 333301
rect 248643 333236 248644 333300
rect 248708 333236 248709 333300
rect 248643 333235 248709 333236
rect 248646 13293 248706 333235
rect 248827 333164 248893 333165
rect 248827 333100 248828 333164
rect 248892 333100 248893 333164
rect 248827 333099 248893 333100
rect 248830 13429 248890 333099
rect 249294 322954 249914 336000
rect 249294 322718 249326 322954
rect 249562 322718 249646 322954
rect 249882 322718 249914 322954
rect 249294 322634 249914 322718
rect 249294 322398 249326 322634
rect 249562 322398 249646 322634
rect 249882 322398 249914 322634
rect 249294 286954 249914 322398
rect 249294 286718 249326 286954
rect 249562 286718 249646 286954
rect 249882 286718 249914 286954
rect 249294 286634 249914 286718
rect 249294 286398 249326 286634
rect 249562 286398 249646 286634
rect 249882 286398 249914 286634
rect 249294 250954 249914 286398
rect 249294 250718 249326 250954
rect 249562 250718 249646 250954
rect 249882 250718 249914 250954
rect 249294 250634 249914 250718
rect 249294 250398 249326 250634
rect 249562 250398 249646 250634
rect 249882 250398 249914 250634
rect 249294 214954 249914 250398
rect 249294 214718 249326 214954
rect 249562 214718 249646 214954
rect 249882 214718 249914 214954
rect 249294 214634 249914 214718
rect 249294 214398 249326 214634
rect 249562 214398 249646 214634
rect 249882 214398 249914 214634
rect 249294 178954 249914 214398
rect 249294 178718 249326 178954
rect 249562 178718 249646 178954
rect 249882 178718 249914 178954
rect 249294 178634 249914 178718
rect 249294 178398 249326 178634
rect 249562 178398 249646 178634
rect 249882 178398 249914 178634
rect 249294 142954 249914 178398
rect 249294 142718 249326 142954
rect 249562 142718 249646 142954
rect 249882 142718 249914 142954
rect 249294 142634 249914 142718
rect 249294 142398 249326 142634
rect 249562 142398 249646 142634
rect 249882 142398 249914 142634
rect 249294 106954 249914 142398
rect 249294 106718 249326 106954
rect 249562 106718 249646 106954
rect 249882 106718 249914 106954
rect 249294 106634 249914 106718
rect 249294 106398 249326 106634
rect 249562 106398 249646 106634
rect 249882 106398 249914 106634
rect 249294 70954 249914 106398
rect 249294 70718 249326 70954
rect 249562 70718 249646 70954
rect 249882 70718 249914 70954
rect 249294 70634 249914 70718
rect 249294 70398 249326 70634
rect 249562 70398 249646 70634
rect 249882 70398 249914 70634
rect 249294 34954 249914 70398
rect 249294 34718 249326 34954
rect 249562 34718 249646 34954
rect 249882 34718 249914 34954
rect 249294 34634 249914 34718
rect 249294 34398 249326 34634
rect 249562 34398 249646 34634
rect 249882 34398 249914 34634
rect 248827 13428 248893 13429
rect 248827 13364 248828 13428
rect 248892 13364 248893 13428
rect 248827 13363 248893 13364
rect 248643 13292 248709 13293
rect 248643 13228 248644 13292
rect 248708 13228 248709 13292
rect 248643 13227 248709 13228
rect 247355 13156 247421 13157
rect 247355 13092 247356 13156
rect 247420 13092 247421 13156
rect 247355 13091 247421 13092
rect 245883 13020 245949 13021
rect 245883 12956 245884 13020
rect 245948 12956 245949 13020
rect 245883 12955 245949 12956
rect 245699 4860 245765 4861
rect 245699 4796 245700 4860
rect 245764 4796 245765 4860
rect 245699 4795 245765 4796
rect 244794 -6342 244826 -6106
rect 245062 -6342 245146 -6106
rect 245382 -6342 245414 -6106
rect 244794 -6426 245414 -6342
rect 244794 -6662 244826 -6426
rect 245062 -6662 245146 -6426
rect 245382 -6662 245414 -6426
rect 244794 -7654 245414 -6662
rect 249294 -7066 249914 34398
rect 250118 13565 250178 337859
rect 250299 337516 250365 337517
rect 250299 337452 250300 337516
rect 250364 337452 250365 337516
rect 250299 337451 250365 337452
rect 250302 177309 250362 337451
rect 251219 333300 251285 333301
rect 251219 333236 251220 333300
rect 251284 333236 251285 333300
rect 251219 333235 251285 333236
rect 250299 177308 250365 177309
rect 250299 177244 250300 177308
rect 250364 177244 250365 177308
rect 250299 177243 250365 177244
rect 250115 13564 250181 13565
rect 250115 13500 250116 13564
rect 250180 13500 250181 13564
rect 250115 13499 250181 13500
rect 251222 10437 251282 333235
rect 251219 10436 251285 10437
rect 251219 10372 251220 10436
rect 251284 10372 251285 10436
rect 251219 10371 251285 10372
rect 251406 10301 251466 337859
rect 251587 337380 251653 337381
rect 251587 337316 251588 337380
rect 251652 337316 251653 337380
rect 251587 337315 251653 337316
rect 251590 14517 251650 337315
rect 251774 80749 251834 337859
rect 252691 337652 252757 337653
rect 252691 337588 252692 337652
rect 252756 337588 252757 337652
rect 252691 337587 252757 337588
rect 252507 334796 252573 334797
rect 252507 334732 252508 334796
rect 252572 334732 252573 334796
rect 252507 334731 252573 334732
rect 251771 80748 251837 80749
rect 251771 80684 251772 80748
rect 251836 80684 251837 80748
rect 251771 80683 251837 80684
rect 251587 14516 251653 14517
rect 251587 14452 251588 14516
rect 251652 14452 251653 14516
rect 251587 14451 251653 14452
rect 251403 10300 251469 10301
rect 251403 10236 251404 10300
rect 251468 10236 251469 10300
rect 251403 10235 251469 10236
rect 252510 4997 252570 334731
rect 252694 7581 252754 337587
rect 252878 327861 252938 337859
rect 254166 336293 254226 337859
rect 254163 336292 254229 336293
rect 254163 336228 254164 336292
rect 254228 336228 254229 336292
rect 254163 336227 254229 336228
rect 252875 327860 252941 327861
rect 252875 327796 252876 327860
rect 252940 327796 252941 327860
rect 252875 327795 252941 327796
rect 253794 327454 254414 336000
rect 253794 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 254414 327454
rect 253794 327134 254414 327218
rect 253794 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 254414 327134
rect 253794 291454 254414 326898
rect 253794 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 254414 291454
rect 253794 291134 254414 291218
rect 253794 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 254414 291134
rect 253794 255454 254414 290898
rect 253794 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 254414 255454
rect 253794 255134 254414 255218
rect 253794 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 254414 255134
rect 253794 219454 254414 254898
rect 253794 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 254414 219454
rect 253794 219134 254414 219218
rect 253794 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 254414 219134
rect 253794 183454 254414 218898
rect 253794 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 254414 183454
rect 253794 183134 254414 183218
rect 253794 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 254414 183134
rect 253794 147454 254414 182898
rect 253794 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 254414 147454
rect 253794 147134 254414 147218
rect 253794 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 254414 147134
rect 253794 111454 254414 146898
rect 253794 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 254414 111454
rect 253794 111134 254414 111218
rect 253794 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 254414 111134
rect 253794 75454 254414 110898
rect 253794 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 254414 75454
rect 253794 75134 254414 75218
rect 253794 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 254414 75134
rect 253794 39454 254414 74898
rect 253794 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 254414 39454
rect 253794 39134 254414 39218
rect 253794 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 254414 39134
rect 252691 7580 252757 7581
rect 252691 7516 252692 7580
rect 252756 7516 252757 7580
rect 252691 7515 252757 7516
rect 252507 4996 252573 4997
rect 252507 4932 252508 4996
rect 252572 4932 252573 4996
rect 252507 4931 252573 4932
rect 249294 -7302 249326 -7066
rect 249562 -7302 249646 -7066
rect 249882 -7302 249914 -7066
rect 249294 -7386 249914 -7302
rect 249294 -7622 249326 -7386
rect 249562 -7622 249646 -7386
rect 249882 -7622 249914 -7386
rect 249294 -7654 249914 -7622
rect 253794 3454 254414 38898
rect 254534 13701 254594 338131
rect 254715 337924 254781 337925
rect 254715 337860 254716 337924
rect 254780 337860 254781 337924
rect 254715 337859 254781 337860
rect 254718 335885 254778 337859
rect 255451 337788 255517 337789
rect 255451 337724 255452 337788
rect 255516 337724 255517 337788
rect 255451 337723 255517 337724
rect 254715 335884 254781 335885
rect 254715 335820 254716 335884
rect 254780 335820 254781 335884
rect 254715 335819 254781 335820
rect 255267 335884 255333 335885
rect 255267 335820 255268 335884
rect 255332 335820 255333 335884
rect 255267 335819 255333 335820
rect 254899 334524 254965 334525
rect 254899 334460 254900 334524
rect 254964 334460 254965 334524
rect 254899 334459 254965 334460
rect 254715 332892 254781 332893
rect 254715 332828 254716 332892
rect 254780 332828 254781 332892
rect 254715 332827 254781 332828
rect 254718 44845 254778 332827
rect 254902 327997 254962 334459
rect 254899 327996 254965 327997
rect 254899 327932 254900 327996
rect 254964 327932 254965 327996
rect 254899 327931 254965 327932
rect 254715 44844 254781 44845
rect 254715 44780 254716 44844
rect 254780 44780 254781 44844
rect 254715 44779 254781 44780
rect 254531 13700 254597 13701
rect 254531 13636 254532 13700
rect 254596 13636 254597 13700
rect 254531 13635 254597 13636
rect 255270 3501 255330 335819
rect 255454 9621 255514 337723
rect 255638 326501 255698 338131
rect 255819 338060 255885 338061
rect 255819 337996 255820 338060
rect 255884 337996 255885 338060
rect 255819 337995 255885 337996
rect 266491 338060 266557 338061
rect 266491 337996 266492 338060
rect 266556 337996 266557 338060
rect 266491 337995 266557 337996
rect 288022 337998 288450 338058
rect 255822 330445 255882 337995
rect 257107 337924 257173 337925
rect 257107 337860 257108 337924
rect 257172 337860 257173 337924
rect 257107 337859 257173 337860
rect 259131 337924 259197 337925
rect 259131 337860 259132 337924
rect 259196 337860 259197 337924
rect 259683 337924 259749 337925
rect 259683 337922 259684 337924
rect 259131 337859 259197 337860
rect 259502 337862 259684 337922
rect 256923 335340 256989 335341
rect 256923 335276 256924 335340
rect 256988 335276 256989 335340
rect 256923 335275 256989 335276
rect 256739 334796 256805 334797
rect 256739 334732 256740 334796
rect 256804 334732 256805 334796
rect 256739 334731 256805 334732
rect 255819 330444 255885 330445
rect 255819 330380 255820 330444
rect 255884 330380 255885 330444
rect 255819 330379 255885 330380
rect 255635 326500 255701 326501
rect 255635 326436 255636 326500
rect 255700 326436 255701 326500
rect 255635 326435 255701 326436
rect 255451 9620 255517 9621
rect 255451 9556 255452 9620
rect 255516 9556 255517 9620
rect 255451 9555 255517 9556
rect 256742 5133 256802 334731
rect 256926 328133 256986 335275
rect 257110 330581 257170 337859
rect 258027 336564 258093 336565
rect 258027 336500 258028 336564
rect 258092 336500 258093 336564
rect 258027 336499 258093 336500
rect 257107 330580 257173 330581
rect 257107 330516 257108 330580
rect 257172 330516 257173 330580
rect 257107 330515 257173 330516
rect 256923 328132 256989 328133
rect 256923 328068 256924 328132
rect 256988 328068 256989 328132
rect 256923 328067 256989 328068
rect 258030 321570 258090 336499
rect 257846 321510 258090 321570
rect 258294 331954 258914 336000
rect 258294 331718 258326 331954
rect 258562 331718 258646 331954
rect 258882 331718 258914 331954
rect 258294 331634 258914 331718
rect 258294 331398 258326 331634
rect 258562 331398 258646 331634
rect 258882 331398 258914 331634
rect 257846 161490 257906 321510
rect 257478 161430 257906 161490
rect 258294 295954 258914 331398
rect 258294 295718 258326 295954
rect 258562 295718 258646 295954
rect 258882 295718 258914 295954
rect 258294 295634 258914 295718
rect 258294 295398 258326 295634
rect 258562 295398 258646 295634
rect 258882 295398 258914 295634
rect 258294 259954 258914 295398
rect 258294 259718 258326 259954
rect 258562 259718 258646 259954
rect 258882 259718 258914 259954
rect 258294 259634 258914 259718
rect 258294 259398 258326 259634
rect 258562 259398 258646 259634
rect 258882 259398 258914 259634
rect 258294 223954 258914 259398
rect 258294 223718 258326 223954
rect 258562 223718 258646 223954
rect 258882 223718 258914 223954
rect 258294 223634 258914 223718
rect 258294 223398 258326 223634
rect 258562 223398 258646 223634
rect 258882 223398 258914 223634
rect 258294 187954 258914 223398
rect 258294 187718 258326 187954
rect 258562 187718 258646 187954
rect 258882 187718 258914 187954
rect 258294 187634 258914 187718
rect 258294 187398 258326 187634
rect 258562 187398 258646 187634
rect 258882 187398 258914 187634
rect 257478 151877 257538 161430
rect 258294 158000 258914 187398
rect 257843 155820 257909 155821
rect 257843 155756 257844 155820
rect 257908 155756 257909 155820
rect 257843 155755 257909 155756
rect 257659 153916 257725 153917
rect 257659 153852 257660 153916
rect 257724 153852 257725 153916
rect 257659 153851 257725 153852
rect 257475 151876 257541 151877
rect 257475 151812 257476 151876
rect 257540 151812 257541 151876
rect 257475 151811 257541 151812
rect 257475 151740 257541 151741
rect 257475 151676 257476 151740
rect 257540 151676 257541 151740
rect 257475 151675 257541 151676
rect 257478 142221 257538 151675
rect 257475 142220 257541 142221
rect 257475 142156 257476 142220
rect 257540 142156 257541 142220
rect 257475 142155 257541 142156
rect 256739 5132 256805 5133
rect 256739 5068 256740 5132
rect 256804 5068 256805 5132
rect 256739 5067 256805 5068
rect 257662 3501 257722 153851
rect 257846 3637 257906 155755
rect 258027 151876 258093 151877
rect 258027 151812 258028 151876
rect 258092 151812 258093 151876
rect 258027 151811 258093 151812
rect 258030 151741 258090 151811
rect 258027 151740 258093 151741
rect 258027 151676 258028 151740
rect 258092 151676 258093 151740
rect 258027 151675 258093 151676
rect 258027 142220 258093 142221
rect 258027 142156 258028 142220
rect 258092 142156 258093 142220
rect 258027 142155 258093 142156
rect 258030 141949 258090 142155
rect 258027 141948 258093 141949
rect 258027 141884 258028 141948
rect 258092 141884 258093 141948
rect 258027 141883 258093 141884
rect 258027 132564 258093 132565
rect 258027 132500 258028 132564
rect 258092 132500 258093 132564
rect 258027 132499 258093 132500
rect 258030 132429 258090 132499
rect 258027 132428 258093 132429
rect 258027 132364 258028 132428
rect 258092 132364 258093 132428
rect 258027 132363 258093 132364
rect 258027 122908 258093 122909
rect 258027 122844 258028 122908
rect 258092 122844 258093 122908
rect 258027 122843 258093 122844
rect 258030 122773 258090 122843
rect 258027 122772 258093 122773
rect 258027 122708 258028 122772
rect 258092 122708 258093 122772
rect 258027 122707 258093 122708
rect 258027 113252 258093 113253
rect 258027 113188 258028 113252
rect 258092 113188 258093 113252
rect 258027 113187 258093 113188
rect 258030 113117 258090 113187
rect 258027 113116 258093 113117
rect 258027 113052 258028 113116
rect 258092 113052 258093 113116
rect 258027 113051 258093 113052
rect 258027 103596 258093 103597
rect 258027 103532 258028 103596
rect 258092 103532 258093 103596
rect 258027 103531 258093 103532
rect 258030 103461 258090 103531
rect 258027 103460 258093 103461
rect 258027 103396 258028 103460
rect 258092 103396 258093 103460
rect 258027 103395 258093 103396
rect 258027 93940 258093 93941
rect 258027 93876 258028 93940
rect 258092 93876 258093 93940
rect 258027 93875 258093 93876
rect 258030 93669 258090 93875
rect 258027 93668 258093 93669
rect 258027 93604 258028 93668
rect 258092 93604 258093 93668
rect 258027 93603 258093 93604
rect 258027 84284 258093 84285
rect 258027 84220 258028 84284
rect 258092 84220 258093 84284
rect 258027 84219 258093 84220
rect 258030 84149 258090 84219
rect 258027 84148 258093 84149
rect 258027 84084 258028 84148
rect 258092 84084 258093 84148
rect 258027 84083 258093 84084
rect 258294 79954 258914 98000
rect 258294 79718 258326 79954
rect 258562 79718 258646 79954
rect 258882 79718 258914 79954
rect 258294 79634 258914 79718
rect 258294 79398 258326 79634
rect 258562 79398 258646 79634
rect 258882 79398 258914 79634
rect 258027 74764 258093 74765
rect 258027 74700 258028 74764
rect 258092 74700 258093 74764
rect 258027 74699 258093 74700
rect 258030 74493 258090 74699
rect 258027 74492 258093 74493
rect 258027 74428 258028 74492
rect 258092 74428 258093 74492
rect 258027 74427 258093 74428
rect 258027 65108 258093 65109
rect 258027 65044 258028 65108
rect 258092 65044 258093 65108
rect 258027 65043 258093 65044
rect 258030 64701 258090 65043
rect 258027 64700 258093 64701
rect 258027 64636 258028 64700
rect 258092 64636 258093 64700
rect 258027 64635 258093 64636
rect 258027 55316 258093 55317
rect 258027 55252 258028 55316
rect 258092 55252 258093 55316
rect 258027 55251 258093 55252
rect 258030 55045 258090 55251
rect 258027 55044 258093 55045
rect 258027 54980 258028 55044
rect 258092 54980 258093 55044
rect 258027 54979 258093 54980
rect 258027 45660 258093 45661
rect 258027 45596 258028 45660
rect 258092 45596 258093 45660
rect 258027 45595 258093 45596
rect 258030 45389 258090 45595
rect 258027 45388 258093 45389
rect 258027 45324 258028 45388
rect 258092 45324 258093 45388
rect 258027 45323 258093 45324
rect 258294 43954 258914 79398
rect 258294 43718 258326 43954
rect 258562 43718 258646 43954
rect 258882 43718 258914 43954
rect 258294 43634 258914 43718
rect 258294 43398 258326 43634
rect 258562 43398 258646 43634
rect 258882 43398 258914 43634
rect 258027 36004 258093 36005
rect 258027 35940 258028 36004
rect 258092 35940 258093 36004
rect 258027 35939 258093 35940
rect 258030 35733 258090 35939
rect 258027 35732 258093 35733
rect 258027 35668 258028 35732
rect 258092 35668 258093 35732
rect 258027 35667 258093 35668
rect 258027 26348 258093 26349
rect 258027 26284 258028 26348
rect 258092 26284 258093 26348
rect 258027 26283 258093 26284
rect 258030 26213 258090 26283
rect 258027 26212 258093 26213
rect 258027 26148 258028 26212
rect 258092 26148 258093 26212
rect 258027 26147 258093 26148
rect 258027 16828 258093 16829
rect 258027 16764 258028 16828
rect 258092 16764 258093 16828
rect 258027 16763 258093 16764
rect 258030 16421 258090 16763
rect 258027 16420 258093 16421
rect 258027 16356 258028 16420
rect 258092 16356 258093 16420
rect 258027 16355 258093 16356
rect 258294 7954 258914 43398
rect 258294 7718 258326 7954
rect 258562 7718 258646 7954
rect 258882 7718 258914 7954
rect 258294 7634 258914 7718
rect 259134 7717 259194 337859
rect 259502 335885 259562 337862
rect 259683 337860 259684 337862
rect 259748 337860 259749 337924
rect 259683 337859 259749 337860
rect 261155 337924 261221 337925
rect 261155 337860 261156 337924
rect 261220 337860 261221 337924
rect 261155 337859 261221 337860
rect 262259 337924 262325 337925
rect 262259 337860 262260 337924
rect 262324 337860 262325 337924
rect 262259 337859 262325 337860
rect 262443 337924 262509 337925
rect 262443 337860 262444 337924
rect 262508 337860 262509 337924
rect 262443 337859 262509 337860
rect 264099 337924 264165 337925
rect 264099 337860 264100 337924
rect 264164 337860 264165 337924
rect 264099 337859 264165 337860
rect 259683 337788 259749 337789
rect 259683 337724 259684 337788
rect 259748 337724 259749 337788
rect 259683 337723 259749 337724
rect 259499 335884 259565 335885
rect 259499 335820 259500 335884
rect 259564 335820 259565 335884
rect 259499 335819 259565 335820
rect 259499 334524 259565 334525
rect 259499 334460 259500 334524
rect 259564 334460 259565 334524
rect 259499 334459 259565 334460
rect 259502 155277 259562 334459
rect 259686 155413 259746 337723
rect 260787 337652 260853 337653
rect 260787 337588 260788 337652
rect 260852 337588 260853 337652
rect 260787 337587 260853 337588
rect 259867 335748 259933 335749
rect 259867 335684 259868 335748
rect 259932 335684 259933 335748
rect 259867 335683 259933 335684
rect 259870 326637 259930 335683
rect 260790 331941 260850 337587
rect 260971 335340 261037 335341
rect 260971 335276 260972 335340
rect 261036 335276 261037 335340
rect 260971 335275 261037 335276
rect 260787 331940 260853 331941
rect 260787 331876 260788 331940
rect 260852 331876 260853 331940
rect 260787 331875 260853 331876
rect 259867 326636 259933 326637
rect 259867 326572 259868 326636
rect 259932 326572 259933 326636
rect 259867 326571 259933 326572
rect 260974 156637 261034 335275
rect 260971 156636 261037 156637
rect 260971 156572 260972 156636
rect 261036 156572 261037 156636
rect 260971 156571 261037 156572
rect 260419 155684 260485 155685
rect 260419 155620 260420 155684
rect 260484 155620 260485 155684
rect 260419 155619 260485 155620
rect 259683 155412 259749 155413
rect 259683 155348 259684 155412
rect 259748 155348 259749 155412
rect 259683 155347 259749 155348
rect 259499 155276 259565 155277
rect 259499 155212 259500 155276
rect 259564 155212 259565 155276
rect 259499 155211 259565 155212
rect 259131 7716 259197 7717
rect 259131 7652 259132 7716
rect 259196 7652 259197 7716
rect 259131 7651 259197 7652
rect 258294 7398 258326 7634
rect 258562 7398 258646 7634
rect 258882 7398 258914 7634
rect 258027 7036 258093 7037
rect 258027 6972 258028 7036
rect 258092 6972 258093 7036
rect 258027 6971 258093 6972
rect 258030 6765 258090 6971
rect 258027 6764 258093 6765
rect 258027 6700 258028 6764
rect 258092 6700 258093 6764
rect 258027 6699 258093 6700
rect 257843 3636 257909 3637
rect 257843 3572 257844 3636
rect 257908 3572 257909 3636
rect 257843 3571 257909 3572
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 255267 3500 255333 3501
rect 255267 3436 255268 3500
rect 255332 3436 255333 3500
rect 255267 3435 255333 3436
rect 257659 3500 257725 3501
rect 257659 3436 257660 3500
rect 257724 3436 257725 3500
rect 257659 3435 257725 3436
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -7654 254414 -902
rect 258294 -1306 258914 7398
rect 260422 3909 260482 155619
rect 261158 155549 261218 337859
rect 262262 157997 262322 337859
rect 262446 335885 262506 337859
rect 263731 337788 263797 337789
rect 263731 337724 263732 337788
rect 263796 337724 263797 337788
rect 263731 337723 263797 337724
rect 262627 336292 262693 336293
rect 262627 336228 262628 336292
rect 262692 336228 262693 336292
rect 262627 336227 262693 336228
rect 262443 335884 262509 335885
rect 262443 335820 262444 335884
rect 262508 335820 262509 335884
rect 262443 335819 262509 335820
rect 262630 160989 262690 336227
rect 262794 300454 263414 336000
rect 263547 331260 263613 331261
rect 263547 331196 263548 331260
rect 263612 331196 263613 331260
rect 263547 331195 263613 331196
rect 263550 331125 263610 331195
rect 263547 331124 263613 331125
rect 263547 331060 263548 331124
rect 263612 331060 263613 331124
rect 263547 331059 263613 331060
rect 263547 321604 263613 321605
rect 263547 321540 263548 321604
rect 263612 321540 263613 321604
rect 263547 321539 263613 321540
rect 262794 300218 262826 300454
rect 263062 300218 263146 300454
rect 263382 300218 263414 300454
rect 262794 300134 263414 300218
rect 262794 299898 262826 300134
rect 263062 299898 263146 300134
rect 263382 299898 263414 300134
rect 262794 264454 263414 299898
rect 262794 264218 262826 264454
rect 263062 264218 263146 264454
rect 263382 264218 263414 264454
rect 262794 264134 263414 264218
rect 262794 263898 262826 264134
rect 263062 263898 263146 264134
rect 263382 263898 263414 264134
rect 262794 228454 263414 263898
rect 262794 228218 262826 228454
rect 263062 228218 263146 228454
rect 263382 228218 263414 228454
rect 262794 228134 263414 228218
rect 262794 227898 262826 228134
rect 263062 227898 263146 228134
rect 263382 227898 263414 228134
rect 262794 192454 263414 227898
rect 262794 192218 262826 192454
rect 263062 192218 263146 192454
rect 263382 192218 263414 192454
rect 262794 192134 263414 192218
rect 262794 191898 262826 192134
rect 263062 191898 263146 192134
rect 263382 191898 263414 192134
rect 262627 160988 262693 160989
rect 262627 160924 262628 160988
rect 262692 160924 262693 160988
rect 262627 160923 262693 160924
rect 262794 158000 263414 191898
rect 263550 158133 263610 321539
rect 263734 159357 263794 337723
rect 263915 336700 263981 336701
rect 263915 336636 263916 336700
rect 263980 336636 263981 336700
rect 263915 336635 263981 336636
rect 263918 328269 263978 336635
rect 264102 331261 264162 337859
rect 265571 337516 265637 337517
rect 265571 337452 265572 337516
rect 265636 337452 265637 337516
rect 265571 337451 265637 337452
rect 265203 335612 265269 335613
rect 265203 335548 265204 335612
rect 265268 335548 265269 335612
rect 265203 335547 265269 335548
rect 265019 335476 265085 335477
rect 265019 335412 265020 335476
rect 265084 335412 265085 335476
rect 265019 335411 265085 335412
rect 264099 331260 264165 331261
rect 264099 331196 264100 331260
rect 264164 331196 264165 331260
rect 264099 331195 264165 331196
rect 263915 328268 263981 328269
rect 263915 328204 263916 328268
rect 263980 328204 263981 328268
rect 263915 328203 263981 328204
rect 263731 159356 263797 159357
rect 263731 159292 263732 159356
rect 263796 159292 263797 159356
rect 263731 159291 263797 159292
rect 265022 158677 265082 335411
rect 265206 159493 265266 335547
rect 265387 335476 265453 335477
rect 265387 335412 265388 335476
rect 265452 335412 265453 335476
rect 265387 335411 265453 335412
rect 265203 159492 265269 159493
rect 265203 159428 265204 159492
rect 265268 159428 265269 159492
rect 265203 159427 265269 159428
rect 265390 158813 265450 335411
rect 265574 326365 265634 337451
rect 266307 336700 266373 336701
rect 266307 336636 266308 336700
rect 266372 336636 266373 336700
rect 266307 336635 266373 336636
rect 265571 326364 265637 326365
rect 265571 326300 265572 326364
rect 265636 326300 265637 326364
rect 265571 326299 265637 326300
rect 265387 158812 265453 158813
rect 265387 158748 265388 158812
rect 265452 158748 265453 158812
rect 265387 158747 265453 158748
rect 265019 158676 265085 158677
rect 265019 158612 265020 158676
rect 265084 158612 265085 158676
rect 265019 158611 265085 158612
rect 263547 158132 263613 158133
rect 263547 158068 263548 158132
rect 263612 158068 263613 158132
rect 263547 158067 263613 158068
rect 262259 157996 262325 157997
rect 262259 157932 262260 157996
rect 262324 157932 262325 157996
rect 262259 157931 262325 157932
rect 261155 155548 261221 155549
rect 261155 155484 261156 155548
rect 261220 155484 261221 155548
rect 261155 155483 261221 155484
rect 260603 155412 260669 155413
rect 260603 155348 260604 155412
rect 260668 155348 260669 155412
rect 260603 155347 260669 155348
rect 260419 3908 260485 3909
rect 260419 3844 260420 3908
rect 260484 3844 260485 3908
rect 260419 3843 260485 3844
rect 260606 3773 260666 155347
rect 266310 155141 266370 336635
rect 266494 158269 266554 337995
rect 270171 337924 270237 337925
rect 270171 337860 270172 337924
rect 270236 337860 270237 337924
rect 270171 337859 270237 337860
rect 272379 337924 272445 337925
rect 272379 337860 272380 337924
rect 272444 337860 272445 337924
rect 272379 337859 272445 337860
rect 274035 337924 274101 337925
rect 274035 337860 274036 337924
rect 274100 337860 274101 337924
rect 274035 337859 274101 337860
rect 274955 337924 275021 337925
rect 274955 337860 274956 337924
rect 275020 337860 275021 337924
rect 274955 337859 275021 337860
rect 275875 337924 275941 337925
rect 275875 337860 275876 337924
rect 275940 337860 275941 337924
rect 275875 337859 275941 337860
rect 276059 337924 276125 337925
rect 276059 337860 276060 337924
rect 276124 337860 276125 337924
rect 276059 337859 276125 337860
rect 278635 337924 278701 337925
rect 278635 337860 278636 337924
rect 278700 337860 278701 337924
rect 278635 337859 278701 337860
rect 279739 337924 279805 337925
rect 279739 337860 279740 337924
rect 279804 337860 279805 337924
rect 279739 337859 279805 337860
rect 280843 337924 280909 337925
rect 280843 337860 280844 337924
rect 280908 337860 280909 337924
rect 280843 337859 280909 337860
rect 282315 337924 282381 337925
rect 282315 337860 282316 337924
rect 282380 337860 282381 337924
rect 282315 337859 282381 337860
rect 284707 337924 284773 337925
rect 284707 337860 284708 337924
rect 284772 337860 284773 337924
rect 284707 337859 284773 337860
rect 286363 337924 286429 337925
rect 286363 337860 286364 337924
rect 286428 337860 286429 337924
rect 286363 337859 286429 337860
rect 267294 304954 267914 336000
rect 268147 335748 268213 335749
rect 268147 335684 268148 335748
rect 268212 335684 268213 335748
rect 268147 335683 268213 335684
rect 267294 304718 267326 304954
rect 267562 304718 267646 304954
rect 267882 304718 267914 304954
rect 267294 304634 267914 304718
rect 267294 304398 267326 304634
rect 267562 304398 267646 304634
rect 267882 304398 267914 304634
rect 267294 268954 267914 304398
rect 267294 268718 267326 268954
rect 267562 268718 267646 268954
rect 267882 268718 267914 268954
rect 267294 268634 267914 268718
rect 267294 268398 267326 268634
rect 267562 268398 267646 268634
rect 267882 268398 267914 268634
rect 267294 232954 267914 268398
rect 267294 232718 267326 232954
rect 267562 232718 267646 232954
rect 267882 232718 267914 232954
rect 267294 232634 267914 232718
rect 267294 232398 267326 232634
rect 267562 232398 267646 232634
rect 267882 232398 267914 232634
rect 267294 196954 267914 232398
rect 267294 196718 267326 196954
rect 267562 196718 267646 196954
rect 267882 196718 267914 196954
rect 267294 196634 267914 196718
rect 267294 196398 267326 196634
rect 267562 196398 267646 196634
rect 267882 196398 267914 196634
rect 267294 160954 267914 196398
rect 267294 160718 267326 160954
rect 267562 160718 267646 160954
rect 267882 160718 267914 160954
rect 267294 160634 267914 160718
rect 267294 160398 267326 160634
rect 267562 160398 267646 160634
rect 267882 160398 267914 160634
rect 266491 158268 266557 158269
rect 266491 158204 266492 158268
rect 266556 158204 266557 158268
rect 266491 158203 266557 158204
rect 267294 158000 267914 160398
rect 266307 155140 266373 155141
rect 266307 155076 266308 155140
rect 266372 155076 266373 155140
rect 266307 155075 266373 155076
rect 268150 153781 268210 335683
rect 268331 335612 268397 335613
rect 268331 335548 268332 335612
rect 268396 335548 268397 335612
rect 268331 335547 268397 335548
rect 268334 155957 268394 335547
rect 268515 335476 268581 335477
rect 268515 335412 268516 335476
rect 268580 335412 268581 335476
rect 268515 335411 268581 335412
rect 269067 335476 269133 335477
rect 269067 335412 269068 335476
rect 269132 335412 269133 335476
rect 269067 335411 269133 335412
rect 268518 161125 268578 335411
rect 268515 161124 268581 161125
rect 268515 161060 268516 161124
rect 268580 161060 268581 161124
rect 268515 161059 268581 161060
rect 268331 155956 268397 155957
rect 268331 155892 268332 155956
rect 268396 155892 268397 155956
rect 268331 155891 268397 155892
rect 269070 153917 269130 335411
rect 270174 158133 270234 337859
rect 270355 337788 270421 337789
rect 270355 337724 270356 337788
rect 270420 337724 270421 337788
rect 270355 337723 270421 337724
rect 270171 158132 270237 158133
rect 270171 158068 270172 158132
rect 270236 158068 270237 158132
rect 270171 158067 270237 158068
rect 270358 155549 270418 337723
rect 272382 336157 272442 337859
rect 272379 336156 272445 336157
rect 272379 336092 272380 336156
rect 272444 336092 272445 336156
rect 272379 336091 272445 336092
rect 271643 335476 271709 335477
rect 271643 335412 271644 335476
rect 271708 335412 271709 335476
rect 271643 335411 271709 335412
rect 271646 158269 271706 335411
rect 271794 309454 272414 336000
rect 274038 320789 274098 337859
rect 274403 337788 274469 337789
rect 274403 337724 274404 337788
rect 274468 337724 274469 337788
rect 274403 337723 274469 337724
rect 274219 333300 274285 333301
rect 274219 333236 274220 333300
rect 274284 333236 274285 333300
rect 274219 333235 274285 333236
rect 274035 320788 274101 320789
rect 274035 320724 274036 320788
rect 274100 320724 274101 320788
rect 274035 320723 274101 320724
rect 271794 309218 271826 309454
rect 272062 309218 272146 309454
rect 272382 309218 272414 309454
rect 271794 309134 272414 309218
rect 271794 308898 271826 309134
rect 272062 308898 272146 309134
rect 272382 308898 272414 309134
rect 271794 273454 272414 308898
rect 271794 273218 271826 273454
rect 272062 273218 272146 273454
rect 272382 273218 272414 273454
rect 271794 273134 272414 273218
rect 271794 272898 271826 273134
rect 272062 272898 272146 273134
rect 272382 272898 272414 273134
rect 271794 237454 272414 272898
rect 271794 237218 271826 237454
rect 272062 237218 272146 237454
rect 272382 237218 272414 237454
rect 271794 237134 272414 237218
rect 271794 236898 271826 237134
rect 272062 236898 272146 237134
rect 272382 236898 272414 237134
rect 271794 201454 272414 236898
rect 271794 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 272414 201454
rect 271794 201134 272414 201218
rect 271794 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 272414 201134
rect 271794 165454 272414 200898
rect 274222 174725 274282 333235
rect 274219 174724 274285 174725
rect 274219 174660 274220 174724
rect 274284 174660 274285 174724
rect 274219 174659 274285 174660
rect 271794 165218 271826 165454
rect 272062 165218 272146 165454
rect 272382 165218 272414 165454
rect 271794 165134 272414 165218
rect 271794 164898 271826 165134
rect 272062 164898 272146 165134
rect 272382 164898 272414 165134
rect 274406 165069 274466 337723
rect 274771 337516 274837 337517
rect 274771 337452 274772 337516
rect 274836 337452 274837 337516
rect 274771 337451 274837 337452
rect 274774 335341 274834 337451
rect 274958 335341 275018 337859
rect 274771 335340 274837 335341
rect 274771 335276 274772 335340
rect 274836 335276 274837 335340
rect 274771 335275 274837 335276
rect 274955 335340 275021 335341
rect 274955 335276 274956 335340
rect 275020 335276 275021 335340
rect 274955 335275 275021 335276
rect 274403 165068 274469 165069
rect 274403 165004 274404 165068
rect 274468 165004 274469 165068
rect 274403 165003 274469 165004
rect 275878 164933 275938 337859
rect 276062 175949 276122 337859
rect 277163 336020 277229 336021
rect 276294 313954 276914 336000
rect 277163 335956 277164 336020
rect 277228 335956 277229 336020
rect 277163 335955 277229 335956
rect 276294 313718 276326 313954
rect 276562 313718 276646 313954
rect 276882 313718 276914 313954
rect 276294 313634 276914 313718
rect 276294 313398 276326 313634
rect 276562 313398 276646 313634
rect 276882 313398 276914 313634
rect 276294 277954 276914 313398
rect 276294 277718 276326 277954
rect 276562 277718 276646 277954
rect 276882 277718 276914 277954
rect 276294 277634 276914 277718
rect 276294 277398 276326 277634
rect 276562 277398 276646 277634
rect 276882 277398 276914 277634
rect 276294 241954 276914 277398
rect 276294 241718 276326 241954
rect 276562 241718 276646 241954
rect 276882 241718 276914 241954
rect 276294 241634 276914 241718
rect 276294 241398 276326 241634
rect 276562 241398 276646 241634
rect 276882 241398 276914 241634
rect 276294 205954 276914 241398
rect 276294 205718 276326 205954
rect 276562 205718 276646 205954
rect 276882 205718 276914 205954
rect 276294 205634 276914 205718
rect 276294 205398 276326 205634
rect 276562 205398 276646 205634
rect 276882 205398 276914 205634
rect 276059 175948 276125 175949
rect 276059 175884 276060 175948
rect 276124 175884 276125 175948
rect 276059 175883 276125 175884
rect 276294 169954 276914 205398
rect 276294 169718 276326 169954
rect 276562 169718 276646 169954
rect 276882 169718 276914 169954
rect 276294 169634 276914 169718
rect 276294 169398 276326 169634
rect 276562 169398 276646 169634
rect 276882 169398 276914 169634
rect 271643 158268 271709 158269
rect 271643 158204 271644 158268
rect 271708 158204 271709 158268
rect 271643 158203 271709 158204
rect 271794 158000 272414 164898
rect 275875 164932 275941 164933
rect 275875 164868 275876 164932
rect 275940 164868 275941 164932
rect 275875 164867 275941 164868
rect 276294 158000 276914 169398
rect 277166 159629 277226 335955
rect 278451 333300 278517 333301
rect 278451 333236 278452 333300
rect 278516 333236 278517 333300
rect 278451 333235 278517 333236
rect 278454 166565 278514 333235
rect 278451 166564 278517 166565
rect 278451 166500 278452 166564
rect 278516 166500 278517 166564
rect 278451 166499 278517 166500
rect 278638 166429 278698 337859
rect 279555 337652 279621 337653
rect 279555 337588 279556 337652
rect 279620 337588 279621 337652
rect 279555 337587 279621 337588
rect 278635 166428 278701 166429
rect 278635 166364 278636 166428
rect 278700 166364 278701 166428
rect 278635 166363 278701 166364
rect 279558 166293 279618 337587
rect 279742 186965 279802 337859
rect 280846 336701 280906 337859
rect 281579 337788 281645 337789
rect 281579 337724 281580 337788
rect 281644 337724 281645 337788
rect 281579 337723 281645 337724
rect 280843 336700 280909 336701
rect 280843 336636 280844 336700
rect 280908 336636 280909 336700
rect 280843 336635 280909 336636
rect 281582 336565 281642 337723
rect 281579 336564 281645 336565
rect 281579 336500 281580 336564
rect 281644 336500 281645 336564
rect 281579 336499 281645 336500
rect 282318 336021 282378 337859
rect 282499 337788 282565 337789
rect 282499 337724 282500 337788
rect 282564 337724 282565 337788
rect 282499 337723 282565 337724
rect 282315 336020 282381 336021
rect 280794 318454 281414 336000
rect 282315 335956 282316 336020
rect 282380 335956 282381 336020
rect 282315 335955 282381 335956
rect 280794 318218 280826 318454
rect 281062 318218 281146 318454
rect 281382 318218 281414 318454
rect 280794 318134 281414 318218
rect 280794 317898 280826 318134
rect 281062 317898 281146 318134
rect 281382 317898 281414 318134
rect 280794 282454 281414 317898
rect 280794 282218 280826 282454
rect 281062 282218 281146 282454
rect 281382 282218 281414 282454
rect 280794 282134 281414 282218
rect 280794 281898 280826 282134
rect 281062 281898 281146 282134
rect 281382 281898 281414 282134
rect 280794 246454 281414 281898
rect 280794 246218 280826 246454
rect 281062 246218 281146 246454
rect 281382 246218 281414 246454
rect 280794 246134 281414 246218
rect 280794 245898 280826 246134
rect 281062 245898 281146 246134
rect 281382 245898 281414 246134
rect 280794 210454 281414 245898
rect 280794 210218 280826 210454
rect 281062 210218 281146 210454
rect 281382 210218 281414 210454
rect 280794 210134 281414 210218
rect 280794 209898 280826 210134
rect 281062 209898 281146 210134
rect 281382 209898 281414 210134
rect 279739 186964 279805 186965
rect 279739 186900 279740 186964
rect 279804 186900 279805 186964
rect 279739 186899 279805 186900
rect 280794 174454 281414 209898
rect 280794 174218 280826 174454
rect 281062 174218 281146 174454
rect 281382 174218 281414 174454
rect 280794 174134 281414 174218
rect 280794 173898 280826 174134
rect 281062 173898 281146 174134
rect 281382 173898 281414 174134
rect 279555 166292 279621 166293
rect 279555 166228 279556 166292
rect 279620 166228 279621 166292
rect 279555 166227 279621 166228
rect 277163 159628 277229 159629
rect 277163 159564 277164 159628
rect 277228 159564 277229 159628
rect 277163 159563 277229 159564
rect 280794 158000 281414 173898
rect 282502 170373 282562 337723
rect 282683 336836 282749 336837
rect 282683 336772 282684 336836
rect 282748 336772 282749 336836
rect 282683 336771 282749 336772
rect 283419 336836 283485 336837
rect 283419 336772 283420 336836
rect 283484 336772 283485 336836
rect 283419 336771 283485 336772
rect 282499 170372 282565 170373
rect 282499 170308 282500 170372
rect 282564 170308 282565 170372
rect 282499 170307 282565 170308
rect 282686 160853 282746 336771
rect 283422 335477 283482 336771
rect 283603 335884 283669 335885
rect 283603 335820 283604 335884
rect 283668 335820 283669 335884
rect 283603 335819 283669 335820
rect 283419 335476 283485 335477
rect 283419 335412 283420 335476
rect 283484 335412 283485 335476
rect 283419 335411 283485 335412
rect 282683 160852 282749 160853
rect 282683 160788 282684 160852
rect 282748 160788 282749 160852
rect 282683 160787 282749 160788
rect 283606 156637 283666 335819
rect 283787 335612 283853 335613
rect 283787 335548 283788 335612
rect 283852 335548 283853 335612
rect 283787 335547 283853 335548
rect 283790 174589 283850 335547
rect 283971 335476 284037 335477
rect 283971 335412 283972 335476
rect 284036 335412 284037 335476
rect 283971 335411 284037 335412
rect 284155 335476 284221 335477
rect 284155 335412 284156 335476
rect 284220 335412 284221 335476
rect 284155 335411 284221 335412
rect 283787 174588 283853 174589
rect 283787 174524 283788 174588
rect 283852 174524 283853 174588
rect 283787 174523 283853 174524
rect 283974 173501 284034 335411
rect 284158 330581 284218 335411
rect 284155 330580 284221 330581
rect 284155 330516 284156 330580
rect 284220 330516 284221 330580
rect 284155 330515 284221 330516
rect 284710 330445 284770 337859
rect 285443 337788 285509 337789
rect 285443 337724 285444 337788
rect 285508 337724 285509 337788
rect 285443 337723 285509 337724
rect 285075 336836 285141 336837
rect 285075 336772 285076 336836
rect 285140 336772 285141 336836
rect 285075 336771 285141 336772
rect 284891 335612 284957 335613
rect 284891 335548 284892 335612
rect 284956 335548 284957 335612
rect 284891 335547 284957 335548
rect 284707 330444 284773 330445
rect 284707 330380 284708 330444
rect 284772 330380 284773 330444
rect 284707 330379 284773 330380
rect 284894 327725 284954 335547
rect 284891 327724 284957 327725
rect 284891 327660 284892 327724
rect 284956 327660 284957 327724
rect 284891 327659 284957 327660
rect 283971 173500 284037 173501
rect 283971 173436 283972 173500
rect 284036 173436 284037 173500
rect 283971 173435 284037 173436
rect 285078 162349 285138 336771
rect 285446 336429 285506 337723
rect 285443 336428 285509 336429
rect 285443 336364 285444 336428
rect 285508 336364 285509 336428
rect 285443 336363 285509 336364
rect 285294 322954 285914 336000
rect 286366 332610 286426 337859
rect 286731 337788 286797 337789
rect 286731 337724 286732 337788
rect 286796 337724 286797 337788
rect 286731 337723 286797 337724
rect 287835 337788 287901 337789
rect 287835 337724 287836 337788
rect 287900 337724 287901 337788
rect 287835 337723 287901 337724
rect 285294 322718 285326 322954
rect 285562 322718 285646 322954
rect 285882 322718 285914 322954
rect 285294 322634 285914 322718
rect 285294 322398 285326 322634
rect 285562 322398 285646 322634
rect 285882 322398 285914 322634
rect 285294 286954 285914 322398
rect 285294 286718 285326 286954
rect 285562 286718 285646 286954
rect 285882 286718 285914 286954
rect 285294 286634 285914 286718
rect 285294 286398 285326 286634
rect 285562 286398 285646 286634
rect 285882 286398 285914 286634
rect 285294 250954 285914 286398
rect 285294 250718 285326 250954
rect 285562 250718 285646 250954
rect 285882 250718 285914 250954
rect 285294 250634 285914 250718
rect 285294 250398 285326 250634
rect 285562 250398 285646 250634
rect 285882 250398 285914 250634
rect 285294 214954 285914 250398
rect 285294 214718 285326 214954
rect 285562 214718 285646 214954
rect 285882 214718 285914 214954
rect 285294 214634 285914 214718
rect 285294 214398 285326 214634
rect 285562 214398 285646 214634
rect 285882 214398 285914 214634
rect 285294 178954 285914 214398
rect 285294 178718 285326 178954
rect 285562 178718 285646 178954
rect 285882 178718 285914 178954
rect 285294 178634 285914 178718
rect 285294 178398 285326 178634
rect 285562 178398 285646 178634
rect 285882 178398 285914 178634
rect 285075 162348 285141 162349
rect 285075 162284 285076 162348
rect 285140 162284 285141 162348
rect 285075 162283 285141 162284
rect 285294 158000 285914 178398
rect 286182 332550 286426 332610
rect 286182 173365 286242 332550
rect 286179 173364 286245 173365
rect 286179 173300 286180 173364
rect 286244 173300 286245 173364
rect 286179 173299 286245 173300
rect 286734 162213 286794 337723
rect 286915 335204 286981 335205
rect 286915 335140 286916 335204
rect 286980 335140 286981 335204
rect 286915 335139 286981 335140
rect 286731 162212 286797 162213
rect 286731 162148 286732 162212
rect 286796 162148 286797 162212
rect 286731 162147 286797 162148
rect 286918 159493 286978 335139
rect 287838 160717 287898 337723
rect 288022 177309 288082 337998
rect 288390 337925 288450 337998
rect 288203 337924 288269 337925
rect 288203 337860 288204 337924
rect 288268 337860 288269 337924
rect 288203 337859 288269 337860
rect 288387 337924 288453 337925
rect 288387 337860 288388 337924
rect 288452 337860 288453 337924
rect 288387 337859 288453 337860
rect 288206 331941 288266 337859
rect 288203 331940 288269 331941
rect 288203 331876 288204 331940
rect 288268 331876 288269 331940
rect 288203 331875 288269 331876
rect 288019 177308 288085 177309
rect 288019 177244 288020 177308
rect 288084 177244 288085 177308
rect 288019 177243 288085 177244
rect 287835 160716 287901 160717
rect 287835 160652 287836 160716
rect 287900 160652 287901 160716
rect 287835 160651 287901 160652
rect 286915 159492 286981 159493
rect 286915 159428 286916 159492
rect 286980 159428 286981 159492
rect 286915 159427 286981 159428
rect 288758 158405 288818 381923
rect 288942 337381 289002 381923
rect 289491 337924 289557 337925
rect 289491 337860 289492 337924
rect 289556 337860 289557 337924
rect 289491 337859 289557 337860
rect 289307 337788 289373 337789
rect 289307 337786 289308 337788
rect 289126 337726 289308 337786
rect 288939 337380 289005 337381
rect 288939 337316 288940 337380
rect 289004 337316 289005 337380
rect 288939 337315 289005 337316
rect 289126 331805 289186 337726
rect 289307 337724 289308 337726
rect 289372 337724 289373 337788
rect 289307 337723 289373 337724
rect 289307 335068 289373 335069
rect 289307 335004 289308 335068
rect 289372 335004 289373 335068
rect 289307 335003 289373 335004
rect 289123 331804 289189 331805
rect 289123 331740 289124 331804
rect 289188 331740 289189 331804
rect 289123 331739 289189 331740
rect 289310 173229 289370 335003
rect 289307 173228 289373 173229
rect 289307 173164 289308 173228
rect 289372 173164 289373 173228
rect 289307 173163 289373 173164
rect 289494 162077 289554 337859
rect 289794 327454 290414 336000
rect 289794 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 290414 327454
rect 289794 327134 290414 327218
rect 289794 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 290414 327134
rect 289794 291454 290414 326898
rect 289794 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 290414 291454
rect 289794 291134 290414 291218
rect 289794 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 290414 291134
rect 289794 255454 290414 290898
rect 289794 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 290414 255454
rect 289794 255134 290414 255218
rect 289794 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 290414 255134
rect 289794 219454 290414 254898
rect 289794 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 290414 219454
rect 289794 219134 290414 219218
rect 289794 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 290414 219134
rect 289794 183454 290414 218898
rect 289794 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 290414 183454
rect 289794 183134 290414 183218
rect 289794 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 290414 183134
rect 289491 162076 289557 162077
rect 289491 162012 289492 162076
rect 289556 162012 289557 162076
rect 289491 162011 289557 162012
rect 288755 158404 288821 158405
rect 288755 158340 288756 158404
rect 288820 158340 288821 158404
rect 288755 158339 288821 158340
rect 289794 158000 290414 182898
rect 290598 158405 290658 382875
rect 290782 338061 290842 384371
rect 291331 383756 291397 383757
rect 291331 383692 291332 383756
rect 291396 383692 291397 383756
rect 291331 383691 291397 383692
rect 290963 382124 291029 382125
rect 290963 382060 290964 382124
rect 291028 382060 291029 382124
rect 290963 382059 291029 382060
rect 290779 338060 290845 338061
rect 290779 337996 290780 338060
rect 290844 337996 290845 338060
rect 290779 337995 290845 337996
rect 290966 161261 291026 382059
rect 291147 381988 291213 381989
rect 291147 381924 291148 381988
rect 291212 381924 291213 381988
rect 291147 381923 291213 381924
rect 290963 161260 291029 161261
rect 290963 161196 290964 161260
rect 291028 161196 291029 161260
rect 290963 161195 291029 161196
rect 291150 158541 291210 381923
rect 291334 333981 291394 383691
rect 293171 382532 293237 382533
rect 293171 382468 293172 382532
rect 293236 382468 293237 382532
rect 293171 382467 293237 382468
rect 291699 381172 291765 381173
rect 291699 381108 291700 381172
rect 291764 381108 291765 381172
rect 291699 381107 291765 381108
rect 291331 333980 291397 333981
rect 291331 333916 291332 333980
rect 291396 333916 291397 333980
rect 291331 333915 291397 333916
rect 291147 158540 291213 158541
rect 291147 158476 291148 158540
rect 291212 158476 291213 158540
rect 291147 158475 291213 158476
rect 290595 158404 290661 158405
rect 290595 158340 290596 158404
rect 290660 158340 290661 158404
rect 290595 158339 290661 158340
rect 291702 157861 291762 381107
rect 293174 158541 293234 382467
rect 293358 180029 293418 384779
rect 294294 384000 294914 403398
rect 298794 706758 299414 711590
rect 298794 706522 298826 706758
rect 299062 706522 299146 706758
rect 299382 706522 299414 706758
rect 298794 706438 299414 706522
rect 298794 706202 298826 706438
rect 299062 706202 299146 706438
rect 299382 706202 299414 706438
rect 298794 696454 299414 706202
rect 298794 696218 298826 696454
rect 299062 696218 299146 696454
rect 299382 696218 299414 696454
rect 298794 696134 299414 696218
rect 298794 695898 298826 696134
rect 299062 695898 299146 696134
rect 299382 695898 299414 696134
rect 298794 660454 299414 695898
rect 298794 660218 298826 660454
rect 299062 660218 299146 660454
rect 299382 660218 299414 660454
rect 298794 660134 299414 660218
rect 298794 659898 298826 660134
rect 299062 659898 299146 660134
rect 299382 659898 299414 660134
rect 298794 624454 299414 659898
rect 298794 624218 298826 624454
rect 299062 624218 299146 624454
rect 299382 624218 299414 624454
rect 298794 624134 299414 624218
rect 298794 623898 298826 624134
rect 299062 623898 299146 624134
rect 299382 623898 299414 624134
rect 298794 588454 299414 623898
rect 298794 588218 298826 588454
rect 299062 588218 299146 588454
rect 299382 588218 299414 588454
rect 298794 588134 299414 588218
rect 298794 587898 298826 588134
rect 299062 587898 299146 588134
rect 299382 587898 299414 588134
rect 298794 552454 299414 587898
rect 298794 552218 298826 552454
rect 299062 552218 299146 552454
rect 299382 552218 299414 552454
rect 298794 552134 299414 552218
rect 298794 551898 298826 552134
rect 299062 551898 299146 552134
rect 299382 551898 299414 552134
rect 298794 516454 299414 551898
rect 298794 516218 298826 516454
rect 299062 516218 299146 516454
rect 299382 516218 299414 516454
rect 298794 516134 299414 516218
rect 298794 515898 298826 516134
rect 299062 515898 299146 516134
rect 299382 515898 299414 516134
rect 298794 480454 299414 515898
rect 298794 480218 298826 480454
rect 299062 480218 299146 480454
rect 299382 480218 299414 480454
rect 298794 480134 299414 480218
rect 298794 479898 298826 480134
rect 299062 479898 299146 480134
rect 299382 479898 299414 480134
rect 298794 444454 299414 479898
rect 298794 444218 298826 444454
rect 299062 444218 299146 444454
rect 299382 444218 299414 444454
rect 298794 444134 299414 444218
rect 298794 443898 298826 444134
rect 299062 443898 299146 444134
rect 299382 443898 299414 444134
rect 298794 408454 299414 443898
rect 298794 408218 298826 408454
rect 299062 408218 299146 408454
rect 299382 408218 299414 408454
rect 298794 408134 299414 408218
rect 298794 407898 298826 408134
rect 299062 407898 299146 408134
rect 299382 407898 299414 408134
rect 296299 384844 296365 384845
rect 296299 384780 296300 384844
rect 296364 384780 296365 384844
rect 296299 384779 296365 384780
rect 295011 384708 295077 384709
rect 295011 384644 295012 384708
rect 295076 384644 295077 384708
rect 295011 384643 295077 384644
rect 293907 381988 293973 381989
rect 293907 381924 293908 381988
rect 293972 381924 293973 381988
rect 293907 381923 293973 381924
rect 293910 194581 293970 381923
rect 294294 331954 294914 336000
rect 294294 331718 294326 331954
rect 294562 331718 294646 331954
rect 294882 331718 294914 331954
rect 294294 331634 294914 331718
rect 294294 331398 294326 331634
rect 294562 331398 294646 331634
rect 294882 331398 294914 331634
rect 294294 295954 294914 331398
rect 294294 295718 294326 295954
rect 294562 295718 294646 295954
rect 294882 295718 294914 295954
rect 294294 295634 294914 295718
rect 294294 295398 294326 295634
rect 294562 295398 294646 295634
rect 294882 295398 294914 295634
rect 294294 259954 294914 295398
rect 294294 259718 294326 259954
rect 294562 259718 294646 259954
rect 294882 259718 294914 259954
rect 294294 259634 294914 259718
rect 294294 259398 294326 259634
rect 294562 259398 294646 259634
rect 294882 259398 294914 259634
rect 294294 223954 294914 259398
rect 294294 223718 294326 223954
rect 294562 223718 294646 223954
rect 294882 223718 294914 223954
rect 294294 223634 294914 223718
rect 294294 223398 294326 223634
rect 294562 223398 294646 223634
rect 294882 223398 294914 223634
rect 293907 194580 293973 194581
rect 293907 194516 293908 194580
rect 293972 194516 293973 194580
rect 293907 194515 293973 194516
rect 294294 187954 294914 223398
rect 294294 187718 294326 187954
rect 294562 187718 294646 187954
rect 294882 187718 294914 187954
rect 294294 187634 294914 187718
rect 294294 187398 294326 187634
rect 294562 187398 294646 187634
rect 294882 187398 294914 187634
rect 293355 180028 293421 180029
rect 293355 179964 293356 180028
rect 293420 179964 293421 180028
rect 293355 179963 293421 179964
rect 293171 158540 293237 158541
rect 293171 158476 293172 158540
rect 293236 158476 293237 158540
rect 293171 158475 293237 158476
rect 294294 158000 294914 187398
rect 295014 170509 295074 384643
rect 296115 382396 296181 382397
rect 296115 382332 296116 382396
rect 296180 382332 296181 382396
rect 296115 382331 296181 382332
rect 295747 381988 295813 381989
rect 295747 381924 295748 381988
rect 295812 381924 295813 381988
rect 295747 381923 295813 381924
rect 295011 170508 295077 170509
rect 295011 170444 295012 170508
rect 295076 170444 295077 170508
rect 295011 170443 295077 170444
rect 295750 158677 295810 381923
rect 296118 374101 296178 382331
rect 296115 374100 296181 374101
rect 296115 374036 296116 374100
rect 296180 374036 296181 374100
rect 296115 374035 296181 374036
rect 296115 373964 296181 373965
rect 296115 373900 296116 373964
rect 296180 373900 296181 373964
rect 296115 373899 296181 373900
rect 296118 364445 296178 373899
rect 296115 364444 296181 364445
rect 296115 364380 296116 364444
rect 296180 364380 296181 364444
rect 296115 364379 296181 364380
rect 296115 364308 296181 364309
rect 296115 364244 296116 364308
rect 296180 364244 296181 364308
rect 296115 364243 296181 364244
rect 296118 354789 296178 364243
rect 296115 354788 296181 354789
rect 296115 354724 296116 354788
rect 296180 354724 296181 354788
rect 296115 354723 296181 354724
rect 296115 354652 296181 354653
rect 296115 354588 296116 354652
rect 296180 354588 296181 354652
rect 296115 354587 296181 354588
rect 296118 345133 296178 354587
rect 296115 345132 296181 345133
rect 296115 345068 296116 345132
rect 296180 345068 296181 345132
rect 296115 345067 296181 345068
rect 296115 344996 296181 344997
rect 296115 344932 296116 344996
rect 296180 344932 296181 344996
rect 296115 344931 296181 344932
rect 296118 335477 296178 344931
rect 296115 335476 296181 335477
rect 296115 335412 296116 335476
rect 296180 335412 296181 335476
rect 296115 335411 296181 335412
rect 296115 161396 296181 161397
rect 296115 161332 296116 161396
rect 296180 161332 296181 161396
rect 296115 161331 296181 161332
rect 295747 158676 295813 158677
rect 295747 158612 295748 158676
rect 295812 158612 295813 158676
rect 295747 158611 295813 158612
rect 291699 157860 291765 157861
rect 291699 157796 291700 157860
rect 291764 157796 291765 157860
rect 291699 157795 291765 157796
rect 283603 156636 283669 156637
rect 283603 156572 283604 156636
rect 283668 156572 283669 156636
rect 283603 156571 283669 156572
rect 296118 155685 296178 161331
rect 296302 159357 296362 384779
rect 298794 384000 299414 407898
rect 303294 707718 303914 711590
rect 303294 707482 303326 707718
rect 303562 707482 303646 707718
rect 303882 707482 303914 707718
rect 303294 707398 303914 707482
rect 303294 707162 303326 707398
rect 303562 707162 303646 707398
rect 303882 707162 303914 707398
rect 303294 700954 303914 707162
rect 303294 700718 303326 700954
rect 303562 700718 303646 700954
rect 303882 700718 303914 700954
rect 303294 700634 303914 700718
rect 303294 700398 303326 700634
rect 303562 700398 303646 700634
rect 303882 700398 303914 700634
rect 303294 664954 303914 700398
rect 303294 664718 303326 664954
rect 303562 664718 303646 664954
rect 303882 664718 303914 664954
rect 303294 664634 303914 664718
rect 303294 664398 303326 664634
rect 303562 664398 303646 664634
rect 303882 664398 303914 664634
rect 303294 628954 303914 664398
rect 303294 628718 303326 628954
rect 303562 628718 303646 628954
rect 303882 628718 303914 628954
rect 303294 628634 303914 628718
rect 303294 628398 303326 628634
rect 303562 628398 303646 628634
rect 303882 628398 303914 628634
rect 303294 592954 303914 628398
rect 303294 592718 303326 592954
rect 303562 592718 303646 592954
rect 303882 592718 303914 592954
rect 303294 592634 303914 592718
rect 303294 592398 303326 592634
rect 303562 592398 303646 592634
rect 303882 592398 303914 592634
rect 303294 556954 303914 592398
rect 303294 556718 303326 556954
rect 303562 556718 303646 556954
rect 303882 556718 303914 556954
rect 303294 556634 303914 556718
rect 303294 556398 303326 556634
rect 303562 556398 303646 556634
rect 303882 556398 303914 556634
rect 303294 520954 303914 556398
rect 303294 520718 303326 520954
rect 303562 520718 303646 520954
rect 303882 520718 303914 520954
rect 303294 520634 303914 520718
rect 303294 520398 303326 520634
rect 303562 520398 303646 520634
rect 303882 520398 303914 520634
rect 303294 484954 303914 520398
rect 303294 484718 303326 484954
rect 303562 484718 303646 484954
rect 303882 484718 303914 484954
rect 303294 484634 303914 484718
rect 303294 484398 303326 484634
rect 303562 484398 303646 484634
rect 303882 484398 303914 484634
rect 303294 448954 303914 484398
rect 303294 448718 303326 448954
rect 303562 448718 303646 448954
rect 303882 448718 303914 448954
rect 303294 448634 303914 448718
rect 303294 448398 303326 448634
rect 303562 448398 303646 448634
rect 303882 448398 303914 448634
rect 303294 412954 303914 448398
rect 303294 412718 303326 412954
rect 303562 412718 303646 412954
rect 303882 412718 303914 412954
rect 303294 412634 303914 412718
rect 303294 412398 303326 412634
rect 303562 412398 303646 412634
rect 303882 412398 303914 412634
rect 296851 383348 296917 383349
rect 296851 383284 296852 383348
rect 296916 383284 296917 383348
rect 296851 383283 296917 383284
rect 296483 381988 296549 381989
rect 296483 381924 296484 381988
rect 296548 381924 296549 381988
rect 296483 381923 296549 381924
rect 296486 161397 296546 381923
rect 296667 374100 296733 374101
rect 296667 374036 296668 374100
rect 296732 374036 296733 374100
rect 296667 374035 296733 374036
rect 296670 373965 296730 374035
rect 296667 373964 296733 373965
rect 296667 373900 296668 373964
rect 296732 373900 296733 373964
rect 296667 373899 296733 373900
rect 296667 364444 296733 364445
rect 296667 364380 296668 364444
rect 296732 364380 296733 364444
rect 296667 364379 296733 364380
rect 296670 364309 296730 364379
rect 296667 364308 296733 364309
rect 296667 364244 296668 364308
rect 296732 364244 296733 364308
rect 296667 364243 296733 364244
rect 296667 354788 296733 354789
rect 296667 354724 296668 354788
rect 296732 354724 296733 354788
rect 296667 354723 296733 354724
rect 296670 354653 296730 354723
rect 296667 354652 296733 354653
rect 296667 354588 296668 354652
rect 296732 354588 296733 354652
rect 296667 354587 296733 354588
rect 296667 345132 296733 345133
rect 296667 345068 296668 345132
rect 296732 345068 296733 345132
rect 296667 345067 296733 345068
rect 296670 344997 296730 345067
rect 296667 344996 296733 344997
rect 296667 344932 296668 344996
rect 296732 344932 296733 344996
rect 296667 344931 296733 344932
rect 296667 335476 296733 335477
rect 296667 335412 296668 335476
rect 296732 335412 296733 335476
rect 296667 335411 296733 335412
rect 296670 335205 296730 335411
rect 296667 335204 296733 335205
rect 296667 335140 296668 335204
rect 296732 335140 296733 335204
rect 296667 335139 296733 335140
rect 296667 325820 296733 325821
rect 296667 325756 296668 325820
rect 296732 325756 296733 325820
rect 296667 325755 296733 325756
rect 296670 325549 296730 325755
rect 296667 325548 296733 325549
rect 296667 325484 296668 325548
rect 296732 325484 296733 325548
rect 296667 325483 296733 325484
rect 296667 316164 296733 316165
rect 296667 316100 296668 316164
rect 296732 316100 296733 316164
rect 296667 316099 296733 316100
rect 296670 316029 296730 316099
rect 296667 316028 296733 316029
rect 296667 315964 296668 316028
rect 296732 315964 296733 316028
rect 296667 315963 296733 315964
rect 296667 306644 296733 306645
rect 296667 306580 296668 306644
rect 296732 306580 296733 306644
rect 296667 306579 296733 306580
rect 296670 306373 296730 306579
rect 296667 306372 296733 306373
rect 296667 306308 296668 306372
rect 296732 306308 296733 306372
rect 296667 306307 296733 306308
rect 296667 296988 296733 296989
rect 296667 296924 296668 296988
rect 296732 296924 296733 296988
rect 296667 296923 296733 296924
rect 296670 296581 296730 296923
rect 296667 296580 296733 296581
rect 296667 296516 296668 296580
rect 296732 296516 296733 296580
rect 296667 296515 296733 296516
rect 296667 287196 296733 287197
rect 296667 287132 296668 287196
rect 296732 287132 296733 287196
rect 296667 287131 296733 287132
rect 296670 286925 296730 287131
rect 296667 286924 296733 286925
rect 296667 286860 296668 286924
rect 296732 286860 296733 286924
rect 296667 286859 296733 286860
rect 296667 277540 296733 277541
rect 296667 277476 296668 277540
rect 296732 277476 296733 277540
rect 296667 277475 296733 277476
rect 296670 277269 296730 277475
rect 296667 277268 296733 277269
rect 296667 277204 296668 277268
rect 296732 277204 296733 277268
rect 296667 277203 296733 277204
rect 296667 267884 296733 267885
rect 296667 267820 296668 267884
rect 296732 267820 296733 267884
rect 296667 267819 296733 267820
rect 296670 267749 296730 267819
rect 296667 267748 296733 267749
rect 296667 267684 296668 267748
rect 296732 267684 296733 267748
rect 296667 267683 296733 267684
rect 296667 248436 296733 248437
rect 296667 248372 296668 248436
rect 296732 248372 296733 248436
rect 296667 248371 296733 248372
rect 296670 248301 296730 248371
rect 296667 248300 296733 248301
rect 296667 248236 296668 248300
rect 296732 248236 296733 248300
rect 296667 248235 296733 248236
rect 296667 238916 296733 238917
rect 296667 238852 296668 238916
rect 296732 238852 296733 238916
rect 296667 238851 296733 238852
rect 296670 238509 296730 238851
rect 296667 238508 296733 238509
rect 296667 238444 296668 238508
rect 296732 238444 296733 238508
rect 296667 238443 296733 238444
rect 296667 229124 296733 229125
rect 296667 229060 296668 229124
rect 296732 229060 296733 229124
rect 296667 229059 296733 229060
rect 296670 228853 296730 229059
rect 296667 228852 296733 228853
rect 296667 228788 296668 228852
rect 296732 228788 296733 228852
rect 296667 228787 296733 228788
rect 296667 219468 296733 219469
rect 296667 219404 296668 219468
rect 296732 219404 296733 219468
rect 296667 219403 296733 219404
rect 296670 219333 296730 219403
rect 296667 219332 296733 219333
rect 296667 219268 296668 219332
rect 296732 219268 296733 219332
rect 296667 219267 296733 219268
rect 296667 209948 296733 209949
rect 296667 209884 296668 209948
rect 296732 209884 296733 209948
rect 296667 209883 296733 209884
rect 296670 209677 296730 209883
rect 296667 209676 296733 209677
rect 296667 209612 296668 209676
rect 296732 209612 296733 209676
rect 296667 209611 296733 209612
rect 296667 200292 296733 200293
rect 296667 200228 296668 200292
rect 296732 200228 296733 200292
rect 296667 200227 296733 200228
rect 296670 200021 296730 200227
rect 296667 200020 296733 200021
rect 296667 199956 296668 200020
rect 296732 199956 296733 200020
rect 296667 199955 296733 199956
rect 296667 190636 296733 190637
rect 296667 190572 296668 190636
rect 296732 190572 296733 190636
rect 296667 190571 296733 190572
rect 296670 190229 296730 190571
rect 296667 190228 296733 190229
rect 296667 190164 296668 190228
rect 296732 190164 296733 190228
rect 296667 190163 296733 190164
rect 296667 180844 296733 180845
rect 296667 180780 296668 180844
rect 296732 180780 296733 180844
rect 296667 180779 296733 180780
rect 296670 180573 296730 180779
rect 296667 180572 296733 180573
rect 296667 180508 296668 180572
rect 296732 180508 296733 180572
rect 296667 180507 296733 180508
rect 296667 171188 296733 171189
rect 296667 171124 296668 171188
rect 296732 171124 296733 171188
rect 296667 171123 296733 171124
rect 296670 171053 296730 171123
rect 296667 171052 296733 171053
rect 296667 170988 296668 171052
rect 296732 170988 296733 171052
rect 296667 170987 296733 170988
rect 296854 163437 296914 383283
rect 298139 382124 298205 382125
rect 298139 382060 298140 382124
rect 298204 382060 298205 382124
rect 298139 382059 298205 382060
rect 298142 332213 298202 382059
rect 303294 376954 303914 412398
rect 303294 376718 303326 376954
rect 303562 376718 303646 376954
rect 303882 376718 303914 376954
rect 303294 376634 303914 376718
rect 303294 376398 303326 376634
rect 303562 376398 303646 376634
rect 303882 376398 303914 376634
rect 303294 340954 303914 376398
rect 303294 340718 303326 340954
rect 303562 340718 303646 340954
rect 303882 340718 303914 340954
rect 303294 340634 303914 340718
rect 303294 340398 303326 340634
rect 303562 340398 303646 340634
rect 303882 340398 303914 340634
rect 298139 332212 298205 332213
rect 298139 332148 298140 332212
rect 298204 332148 298205 332212
rect 298139 332147 298205 332148
rect 298794 300454 299414 336000
rect 298794 300218 298826 300454
rect 299062 300218 299146 300454
rect 299382 300218 299414 300454
rect 298794 300134 299414 300218
rect 298794 299898 298826 300134
rect 299062 299898 299146 300134
rect 299382 299898 299414 300134
rect 298794 264454 299414 299898
rect 298794 264218 298826 264454
rect 299062 264218 299146 264454
rect 299382 264218 299414 264454
rect 298794 264134 299414 264218
rect 298794 263898 298826 264134
rect 299062 263898 299146 264134
rect 299382 263898 299414 264134
rect 298794 228454 299414 263898
rect 298794 228218 298826 228454
rect 299062 228218 299146 228454
rect 299382 228218 299414 228454
rect 298794 228134 299414 228218
rect 298794 227898 298826 228134
rect 299062 227898 299146 228134
rect 299382 227898 299414 228134
rect 298794 192454 299414 227898
rect 298794 192218 298826 192454
rect 299062 192218 299146 192454
rect 299382 192218 299414 192454
rect 298794 192134 299414 192218
rect 298794 191898 298826 192134
rect 299062 191898 299146 192134
rect 299382 191898 299414 192134
rect 296851 163436 296917 163437
rect 296851 163372 296852 163436
rect 296916 163372 296917 163436
rect 296851 163371 296917 163372
rect 296851 161532 296917 161533
rect 296851 161468 296852 161532
rect 296916 161468 296917 161532
rect 296851 161467 296917 161468
rect 296483 161396 296549 161397
rect 296483 161332 296484 161396
rect 296548 161332 296549 161396
rect 296483 161331 296549 161332
rect 296854 160850 296914 161467
rect 296486 160790 296914 160850
rect 296299 159356 296365 159357
rect 296299 159292 296300 159356
rect 296364 159292 296365 159356
rect 296299 159291 296365 159292
rect 296486 158810 296546 160790
rect 296486 158750 296730 158810
rect 296670 158677 296730 158750
rect 296667 158676 296733 158677
rect 296667 158612 296668 158676
rect 296732 158612 296733 158676
rect 296667 158611 296733 158612
rect 298794 158000 299414 191898
rect 303294 304954 303914 340398
rect 303294 304718 303326 304954
rect 303562 304718 303646 304954
rect 303882 304718 303914 304954
rect 303294 304634 303914 304718
rect 303294 304398 303326 304634
rect 303562 304398 303646 304634
rect 303882 304398 303914 304634
rect 303294 268954 303914 304398
rect 303294 268718 303326 268954
rect 303562 268718 303646 268954
rect 303882 268718 303914 268954
rect 303294 268634 303914 268718
rect 303294 268398 303326 268634
rect 303562 268398 303646 268634
rect 303882 268398 303914 268634
rect 303294 232954 303914 268398
rect 303294 232718 303326 232954
rect 303562 232718 303646 232954
rect 303882 232718 303914 232954
rect 303294 232634 303914 232718
rect 303294 232398 303326 232634
rect 303562 232398 303646 232634
rect 303882 232398 303914 232634
rect 303294 196954 303914 232398
rect 303294 196718 303326 196954
rect 303562 196718 303646 196954
rect 303882 196718 303914 196954
rect 303294 196634 303914 196718
rect 303294 196398 303326 196634
rect 303562 196398 303646 196634
rect 303882 196398 303914 196634
rect 303294 160954 303914 196398
rect 303294 160718 303326 160954
rect 303562 160718 303646 160954
rect 303882 160718 303914 160954
rect 303294 160634 303914 160718
rect 303294 160398 303326 160634
rect 303562 160398 303646 160634
rect 303882 160398 303914 160634
rect 303294 158000 303914 160398
rect 307794 708678 308414 711590
rect 307794 708442 307826 708678
rect 308062 708442 308146 708678
rect 308382 708442 308414 708678
rect 307794 708358 308414 708442
rect 307794 708122 307826 708358
rect 308062 708122 308146 708358
rect 308382 708122 308414 708358
rect 307794 669454 308414 708122
rect 307794 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 308414 669454
rect 307794 669134 308414 669218
rect 307794 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 308414 669134
rect 307794 633454 308414 668898
rect 307794 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 308414 633454
rect 307794 633134 308414 633218
rect 307794 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 308414 633134
rect 307794 597454 308414 632898
rect 307794 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 308414 597454
rect 307794 597134 308414 597218
rect 307794 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 308414 597134
rect 307794 561454 308414 596898
rect 307794 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 308414 561454
rect 307794 561134 308414 561218
rect 307794 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 308414 561134
rect 307794 525454 308414 560898
rect 307794 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 308414 525454
rect 307794 525134 308414 525218
rect 307794 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 308414 525134
rect 307794 489454 308414 524898
rect 307794 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 308414 489454
rect 307794 489134 308414 489218
rect 307794 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 308414 489134
rect 307794 453454 308414 488898
rect 307794 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 308414 453454
rect 307794 453134 308414 453218
rect 307794 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 308414 453134
rect 307794 417454 308414 452898
rect 307794 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 308414 417454
rect 307794 417134 308414 417218
rect 307794 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 308414 417134
rect 307794 381454 308414 416898
rect 307794 381218 307826 381454
rect 308062 381218 308146 381454
rect 308382 381218 308414 381454
rect 307794 381134 308414 381218
rect 307794 380898 307826 381134
rect 308062 380898 308146 381134
rect 308382 380898 308414 381134
rect 307794 345454 308414 380898
rect 307794 345218 307826 345454
rect 308062 345218 308146 345454
rect 308382 345218 308414 345454
rect 307794 345134 308414 345218
rect 307794 344898 307826 345134
rect 308062 344898 308146 345134
rect 308382 344898 308414 345134
rect 307794 309454 308414 344898
rect 307794 309218 307826 309454
rect 308062 309218 308146 309454
rect 308382 309218 308414 309454
rect 307794 309134 308414 309218
rect 307794 308898 307826 309134
rect 308062 308898 308146 309134
rect 308382 308898 308414 309134
rect 307794 273454 308414 308898
rect 307794 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 308414 273454
rect 307794 273134 308414 273218
rect 307794 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 308414 273134
rect 307794 237454 308414 272898
rect 307794 237218 307826 237454
rect 308062 237218 308146 237454
rect 308382 237218 308414 237454
rect 307794 237134 308414 237218
rect 307794 236898 307826 237134
rect 308062 236898 308146 237134
rect 308382 236898 308414 237134
rect 307794 201454 308414 236898
rect 307794 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 308414 201454
rect 307794 201134 308414 201218
rect 307794 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 308414 201134
rect 307794 165454 308414 200898
rect 307794 165218 307826 165454
rect 308062 165218 308146 165454
rect 308382 165218 308414 165454
rect 307794 165134 308414 165218
rect 307794 164898 307826 165134
rect 308062 164898 308146 165134
rect 308382 164898 308414 165134
rect 307794 158000 308414 164898
rect 312294 709638 312914 711590
rect 312294 709402 312326 709638
rect 312562 709402 312646 709638
rect 312882 709402 312914 709638
rect 312294 709318 312914 709402
rect 312294 709082 312326 709318
rect 312562 709082 312646 709318
rect 312882 709082 312914 709318
rect 312294 673954 312914 709082
rect 312294 673718 312326 673954
rect 312562 673718 312646 673954
rect 312882 673718 312914 673954
rect 312294 673634 312914 673718
rect 312294 673398 312326 673634
rect 312562 673398 312646 673634
rect 312882 673398 312914 673634
rect 312294 637954 312914 673398
rect 312294 637718 312326 637954
rect 312562 637718 312646 637954
rect 312882 637718 312914 637954
rect 312294 637634 312914 637718
rect 312294 637398 312326 637634
rect 312562 637398 312646 637634
rect 312882 637398 312914 637634
rect 312294 601954 312914 637398
rect 312294 601718 312326 601954
rect 312562 601718 312646 601954
rect 312882 601718 312914 601954
rect 312294 601634 312914 601718
rect 312294 601398 312326 601634
rect 312562 601398 312646 601634
rect 312882 601398 312914 601634
rect 312294 565954 312914 601398
rect 312294 565718 312326 565954
rect 312562 565718 312646 565954
rect 312882 565718 312914 565954
rect 312294 565634 312914 565718
rect 312294 565398 312326 565634
rect 312562 565398 312646 565634
rect 312882 565398 312914 565634
rect 312294 529954 312914 565398
rect 312294 529718 312326 529954
rect 312562 529718 312646 529954
rect 312882 529718 312914 529954
rect 312294 529634 312914 529718
rect 312294 529398 312326 529634
rect 312562 529398 312646 529634
rect 312882 529398 312914 529634
rect 312294 493954 312914 529398
rect 312294 493718 312326 493954
rect 312562 493718 312646 493954
rect 312882 493718 312914 493954
rect 312294 493634 312914 493718
rect 312294 493398 312326 493634
rect 312562 493398 312646 493634
rect 312882 493398 312914 493634
rect 312294 457954 312914 493398
rect 312294 457718 312326 457954
rect 312562 457718 312646 457954
rect 312882 457718 312914 457954
rect 312294 457634 312914 457718
rect 312294 457398 312326 457634
rect 312562 457398 312646 457634
rect 312882 457398 312914 457634
rect 312294 421954 312914 457398
rect 312294 421718 312326 421954
rect 312562 421718 312646 421954
rect 312882 421718 312914 421954
rect 312294 421634 312914 421718
rect 312294 421398 312326 421634
rect 312562 421398 312646 421634
rect 312882 421398 312914 421634
rect 312294 385954 312914 421398
rect 312294 385718 312326 385954
rect 312562 385718 312646 385954
rect 312882 385718 312914 385954
rect 312294 385634 312914 385718
rect 312294 385398 312326 385634
rect 312562 385398 312646 385634
rect 312882 385398 312914 385634
rect 312294 349954 312914 385398
rect 312294 349718 312326 349954
rect 312562 349718 312646 349954
rect 312882 349718 312914 349954
rect 312294 349634 312914 349718
rect 312294 349398 312326 349634
rect 312562 349398 312646 349634
rect 312882 349398 312914 349634
rect 312294 313954 312914 349398
rect 312294 313718 312326 313954
rect 312562 313718 312646 313954
rect 312882 313718 312914 313954
rect 312294 313634 312914 313718
rect 312294 313398 312326 313634
rect 312562 313398 312646 313634
rect 312882 313398 312914 313634
rect 312294 277954 312914 313398
rect 312294 277718 312326 277954
rect 312562 277718 312646 277954
rect 312882 277718 312914 277954
rect 312294 277634 312914 277718
rect 312294 277398 312326 277634
rect 312562 277398 312646 277634
rect 312882 277398 312914 277634
rect 312294 241954 312914 277398
rect 312294 241718 312326 241954
rect 312562 241718 312646 241954
rect 312882 241718 312914 241954
rect 312294 241634 312914 241718
rect 312294 241398 312326 241634
rect 312562 241398 312646 241634
rect 312882 241398 312914 241634
rect 312294 205954 312914 241398
rect 312294 205718 312326 205954
rect 312562 205718 312646 205954
rect 312882 205718 312914 205954
rect 312294 205634 312914 205718
rect 312294 205398 312326 205634
rect 312562 205398 312646 205634
rect 312882 205398 312914 205634
rect 312294 169954 312914 205398
rect 312294 169718 312326 169954
rect 312562 169718 312646 169954
rect 312882 169718 312914 169954
rect 312294 169634 312914 169718
rect 312294 169398 312326 169634
rect 312562 169398 312646 169634
rect 312882 169398 312914 169634
rect 312294 158000 312914 169398
rect 316794 710598 317414 711590
rect 316794 710362 316826 710598
rect 317062 710362 317146 710598
rect 317382 710362 317414 710598
rect 316794 710278 317414 710362
rect 316794 710042 316826 710278
rect 317062 710042 317146 710278
rect 317382 710042 317414 710278
rect 316794 678454 317414 710042
rect 316794 678218 316826 678454
rect 317062 678218 317146 678454
rect 317382 678218 317414 678454
rect 316794 678134 317414 678218
rect 316794 677898 316826 678134
rect 317062 677898 317146 678134
rect 317382 677898 317414 678134
rect 316794 642454 317414 677898
rect 316794 642218 316826 642454
rect 317062 642218 317146 642454
rect 317382 642218 317414 642454
rect 316794 642134 317414 642218
rect 316794 641898 316826 642134
rect 317062 641898 317146 642134
rect 317382 641898 317414 642134
rect 316794 606454 317414 641898
rect 316794 606218 316826 606454
rect 317062 606218 317146 606454
rect 317382 606218 317414 606454
rect 316794 606134 317414 606218
rect 316794 605898 316826 606134
rect 317062 605898 317146 606134
rect 317382 605898 317414 606134
rect 316794 570454 317414 605898
rect 316794 570218 316826 570454
rect 317062 570218 317146 570454
rect 317382 570218 317414 570454
rect 316794 570134 317414 570218
rect 316794 569898 316826 570134
rect 317062 569898 317146 570134
rect 317382 569898 317414 570134
rect 316794 534454 317414 569898
rect 316794 534218 316826 534454
rect 317062 534218 317146 534454
rect 317382 534218 317414 534454
rect 316794 534134 317414 534218
rect 316794 533898 316826 534134
rect 317062 533898 317146 534134
rect 317382 533898 317414 534134
rect 316794 498454 317414 533898
rect 316794 498218 316826 498454
rect 317062 498218 317146 498454
rect 317382 498218 317414 498454
rect 316794 498134 317414 498218
rect 316794 497898 316826 498134
rect 317062 497898 317146 498134
rect 317382 497898 317414 498134
rect 316794 462454 317414 497898
rect 316794 462218 316826 462454
rect 317062 462218 317146 462454
rect 317382 462218 317414 462454
rect 316794 462134 317414 462218
rect 316794 461898 316826 462134
rect 317062 461898 317146 462134
rect 317382 461898 317414 462134
rect 316794 426454 317414 461898
rect 316794 426218 316826 426454
rect 317062 426218 317146 426454
rect 317382 426218 317414 426454
rect 316794 426134 317414 426218
rect 316794 425898 316826 426134
rect 317062 425898 317146 426134
rect 317382 425898 317414 426134
rect 316794 390454 317414 425898
rect 316794 390218 316826 390454
rect 317062 390218 317146 390454
rect 317382 390218 317414 390454
rect 316794 390134 317414 390218
rect 316794 389898 316826 390134
rect 317062 389898 317146 390134
rect 317382 389898 317414 390134
rect 316794 354454 317414 389898
rect 316794 354218 316826 354454
rect 317062 354218 317146 354454
rect 317382 354218 317414 354454
rect 316794 354134 317414 354218
rect 316794 353898 316826 354134
rect 317062 353898 317146 354134
rect 317382 353898 317414 354134
rect 316794 318454 317414 353898
rect 316794 318218 316826 318454
rect 317062 318218 317146 318454
rect 317382 318218 317414 318454
rect 316794 318134 317414 318218
rect 316794 317898 316826 318134
rect 317062 317898 317146 318134
rect 317382 317898 317414 318134
rect 316794 282454 317414 317898
rect 316794 282218 316826 282454
rect 317062 282218 317146 282454
rect 317382 282218 317414 282454
rect 316794 282134 317414 282218
rect 316794 281898 316826 282134
rect 317062 281898 317146 282134
rect 317382 281898 317414 282134
rect 316794 246454 317414 281898
rect 316794 246218 316826 246454
rect 317062 246218 317146 246454
rect 317382 246218 317414 246454
rect 316794 246134 317414 246218
rect 316794 245898 316826 246134
rect 317062 245898 317146 246134
rect 317382 245898 317414 246134
rect 316794 210454 317414 245898
rect 316794 210218 316826 210454
rect 317062 210218 317146 210454
rect 317382 210218 317414 210454
rect 316794 210134 317414 210218
rect 316794 209898 316826 210134
rect 317062 209898 317146 210134
rect 317382 209898 317414 210134
rect 316794 174454 317414 209898
rect 316794 174218 316826 174454
rect 317062 174218 317146 174454
rect 317382 174218 317414 174454
rect 316794 174134 317414 174218
rect 316794 173898 316826 174134
rect 317062 173898 317146 174134
rect 317382 173898 317414 174134
rect 316794 158000 317414 173898
rect 321294 711558 321914 711590
rect 321294 711322 321326 711558
rect 321562 711322 321646 711558
rect 321882 711322 321914 711558
rect 321294 711238 321914 711322
rect 321294 711002 321326 711238
rect 321562 711002 321646 711238
rect 321882 711002 321914 711238
rect 321294 682954 321914 711002
rect 321294 682718 321326 682954
rect 321562 682718 321646 682954
rect 321882 682718 321914 682954
rect 321294 682634 321914 682718
rect 321294 682398 321326 682634
rect 321562 682398 321646 682634
rect 321882 682398 321914 682634
rect 321294 646954 321914 682398
rect 321294 646718 321326 646954
rect 321562 646718 321646 646954
rect 321882 646718 321914 646954
rect 321294 646634 321914 646718
rect 321294 646398 321326 646634
rect 321562 646398 321646 646634
rect 321882 646398 321914 646634
rect 321294 610954 321914 646398
rect 321294 610718 321326 610954
rect 321562 610718 321646 610954
rect 321882 610718 321914 610954
rect 321294 610634 321914 610718
rect 321294 610398 321326 610634
rect 321562 610398 321646 610634
rect 321882 610398 321914 610634
rect 321294 574954 321914 610398
rect 321294 574718 321326 574954
rect 321562 574718 321646 574954
rect 321882 574718 321914 574954
rect 321294 574634 321914 574718
rect 321294 574398 321326 574634
rect 321562 574398 321646 574634
rect 321882 574398 321914 574634
rect 321294 538954 321914 574398
rect 321294 538718 321326 538954
rect 321562 538718 321646 538954
rect 321882 538718 321914 538954
rect 321294 538634 321914 538718
rect 321294 538398 321326 538634
rect 321562 538398 321646 538634
rect 321882 538398 321914 538634
rect 321294 502954 321914 538398
rect 321294 502718 321326 502954
rect 321562 502718 321646 502954
rect 321882 502718 321914 502954
rect 321294 502634 321914 502718
rect 321294 502398 321326 502634
rect 321562 502398 321646 502634
rect 321882 502398 321914 502634
rect 321294 466954 321914 502398
rect 321294 466718 321326 466954
rect 321562 466718 321646 466954
rect 321882 466718 321914 466954
rect 321294 466634 321914 466718
rect 321294 466398 321326 466634
rect 321562 466398 321646 466634
rect 321882 466398 321914 466634
rect 321294 430954 321914 466398
rect 321294 430718 321326 430954
rect 321562 430718 321646 430954
rect 321882 430718 321914 430954
rect 321294 430634 321914 430718
rect 321294 430398 321326 430634
rect 321562 430398 321646 430634
rect 321882 430398 321914 430634
rect 321294 394954 321914 430398
rect 321294 394718 321326 394954
rect 321562 394718 321646 394954
rect 321882 394718 321914 394954
rect 321294 394634 321914 394718
rect 321294 394398 321326 394634
rect 321562 394398 321646 394634
rect 321882 394398 321914 394634
rect 321294 358954 321914 394398
rect 321294 358718 321326 358954
rect 321562 358718 321646 358954
rect 321882 358718 321914 358954
rect 321294 358634 321914 358718
rect 321294 358398 321326 358634
rect 321562 358398 321646 358634
rect 321882 358398 321914 358634
rect 321294 322954 321914 358398
rect 321294 322718 321326 322954
rect 321562 322718 321646 322954
rect 321882 322718 321914 322954
rect 321294 322634 321914 322718
rect 321294 322398 321326 322634
rect 321562 322398 321646 322634
rect 321882 322398 321914 322634
rect 321294 286954 321914 322398
rect 321294 286718 321326 286954
rect 321562 286718 321646 286954
rect 321882 286718 321914 286954
rect 321294 286634 321914 286718
rect 321294 286398 321326 286634
rect 321562 286398 321646 286634
rect 321882 286398 321914 286634
rect 321294 250954 321914 286398
rect 321294 250718 321326 250954
rect 321562 250718 321646 250954
rect 321882 250718 321914 250954
rect 321294 250634 321914 250718
rect 321294 250398 321326 250634
rect 321562 250398 321646 250634
rect 321882 250398 321914 250634
rect 321294 214954 321914 250398
rect 321294 214718 321326 214954
rect 321562 214718 321646 214954
rect 321882 214718 321914 214954
rect 321294 214634 321914 214718
rect 321294 214398 321326 214634
rect 321562 214398 321646 214634
rect 321882 214398 321914 214634
rect 321294 178954 321914 214398
rect 321294 178718 321326 178954
rect 321562 178718 321646 178954
rect 321882 178718 321914 178954
rect 321294 178634 321914 178718
rect 321294 178398 321326 178634
rect 321562 178398 321646 178634
rect 321882 178398 321914 178634
rect 321294 158000 321914 178398
rect 325794 704838 326414 711590
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 687454 326414 704282
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 651454 326414 686898
rect 325794 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 326414 651454
rect 325794 651134 326414 651218
rect 325794 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 326414 651134
rect 325794 615454 326414 650898
rect 325794 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 326414 615454
rect 325794 615134 326414 615218
rect 325794 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 326414 615134
rect 325794 579454 326414 614898
rect 325794 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 326414 579454
rect 325794 579134 326414 579218
rect 325794 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 326414 579134
rect 325794 543454 326414 578898
rect 325794 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 326414 543454
rect 325794 543134 326414 543218
rect 325794 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 326414 543134
rect 325794 507454 326414 542898
rect 325794 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 326414 507454
rect 325794 507134 326414 507218
rect 325794 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 326414 507134
rect 325794 471454 326414 506898
rect 325794 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 326414 471454
rect 325794 471134 326414 471218
rect 325794 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 326414 471134
rect 325794 435454 326414 470898
rect 325794 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 326414 435454
rect 325794 435134 326414 435218
rect 325794 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 326414 435134
rect 325794 399454 326414 434898
rect 325794 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 326414 399454
rect 325794 399134 326414 399218
rect 325794 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 326414 399134
rect 325794 363454 326414 398898
rect 325794 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 326414 363454
rect 325794 363134 326414 363218
rect 325794 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 326414 363134
rect 325794 327454 326414 362898
rect 325794 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 326414 327454
rect 325794 327134 326414 327218
rect 325794 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 326414 327134
rect 325794 291454 326414 326898
rect 325794 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 326414 291454
rect 325794 291134 326414 291218
rect 325794 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 326414 291134
rect 325794 255454 326414 290898
rect 325794 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 326414 255454
rect 325794 255134 326414 255218
rect 325794 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 326414 255134
rect 325794 219454 326414 254898
rect 325794 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 326414 219454
rect 325794 219134 326414 219218
rect 325794 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 326414 219134
rect 325794 183454 326414 218898
rect 325794 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 326414 183454
rect 325794 183134 326414 183218
rect 325794 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 326414 183134
rect 325794 158000 326414 182898
rect 330294 705798 330914 711590
rect 330294 705562 330326 705798
rect 330562 705562 330646 705798
rect 330882 705562 330914 705798
rect 330294 705478 330914 705562
rect 330294 705242 330326 705478
rect 330562 705242 330646 705478
rect 330882 705242 330914 705478
rect 330294 691954 330914 705242
rect 330294 691718 330326 691954
rect 330562 691718 330646 691954
rect 330882 691718 330914 691954
rect 330294 691634 330914 691718
rect 330294 691398 330326 691634
rect 330562 691398 330646 691634
rect 330882 691398 330914 691634
rect 330294 655954 330914 691398
rect 330294 655718 330326 655954
rect 330562 655718 330646 655954
rect 330882 655718 330914 655954
rect 330294 655634 330914 655718
rect 330294 655398 330326 655634
rect 330562 655398 330646 655634
rect 330882 655398 330914 655634
rect 330294 619954 330914 655398
rect 330294 619718 330326 619954
rect 330562 619718 330646 619954
rect 330882 619718 330914 619954
rect 330294 619634 330914 619718
rect 330294 619398 330326 619634
rect 330562 619398 330646 619634
rect 330882 619398 330914 619634
rect 330294 583954 330914 619398
rect 330294 583718 330326 583954
rect 330562 583718 330646 583954
rect 330882 583718 330914 583954
rect 330294 583634 330914 583718
rect 330294 583398 330326 583634
rect 330562 583398 330646 583634
rect 330882 583398 330914 583634
rect 330294 547954 330914 583398
rect 330294 547718 330326 547954
rect 330562 547718 330646 547954
rect 330882 547718 330914 547954
rect 330294 547634 330914 547718
rect 330294 547398 330326 547634
rect 330562 547398 330646 547634
rect 330882 547398 330914 547634
rect 330294 511954 330914 547398
rect 330294 511718 330326 511954
rect 330562 511718 330646 511954
rect 330882 511718 330914 511954
rect 330294 511634 330914 511718
rect 330294 511398 330326 511634
rect 330562 511398 330646 511634
rect 330882 511398 330914 511634
rect 330294 475954 330914 511398
rect 330294 475718 330326 475954
rect 330562 475718 330646 475954
rect 330882 475718 330914 475954
rect 330294 475634 330914 475718
rect 330294 475398 330326 475634
rect 330562 475398 330646 475634
rect 330882 475398 330914 475634
rect 330294 439954 330914 475398
rect 330294 439718 330326 439954
rect 330562 439718 330646 439954
rect 330882 439718 330914 439954
rect 330294 439634 330914 439718
rect 330294 439398 330326 439634
rect 330562 439398 330646 439634
rect 330882 439398 330914 439634
rect 330294 403954 330914 439398
rect 330294 403718 330326 403954
rect 330562 403718 330646 403954
rect 330882 403718 330914 403954
rect 330294 403634 330914 403718
rect 330294 403398 330326 403634
rect 330562 403398 330646 403634
rect 330882 403398 330914 403634
rect 330294 367954 330914 403398
rect 330294 367718 330326 367954
rect 330562 367718 330646 367954
rect 330882 367718 330914 367954
rect 330294 367634 330914 367718
rect 330294 367398 330326 367634
rect 330562 367398 330646 367634
rect 330882 367398 330914 367634
rect 330294 331954 330914 367398
rect 330294 331718 330326 331954
rect 330562 331718 330646 331954
rect 330882 331718 330914 331954
rect 330294 331634 330914 331718
rect 330294 331398 330326 331634
rect 330562 331398 330646 331634
rect 330882 331398 330914 331634
rect 330294 295954 330914 331398
rect 330294 295718 330326 295954
rect 330562 295718 330646 295954
rect 330882 295718 330914 295954
rect 330294 295634 330914 295718
rect 330294 295398 330326 295634
rect 330562 295398 330646 295634
rect 330882 295398 330914 295634
rect 330294 259954 330914 295398
rect 330294 259718 330326 259954
rect 330562 259718 330646 259954
rect 330882 259718 330914 259954
rect 330294 259634 330914 259718
rect 330294 259398 330326 259634
rect 330562 259398 330646 259634
rect 330882 259398 330914 259634
rect 330294 223954 330914 259398
rect 330294 223718 330326 223954
rect 330562 223718 330646 223954
rect 330882 223718 330914 223954
rect 330294 223634 330914 223718
rect 330294 223398 330326 223634
rect 330562 223398 330646 223634
rect 330882 223398 330914 223634
rect 330294 187954 330914 223398
rect 330294 187718 330326 187954
rect 330562 187718 330646 187954
rect 330882 187718 330914 187954
rect 330294 187634 330914 187718
rect 330294 187398 330326 187634
rect 330562 187398 330646 187634
rect 330882 187398 330914 187634
rect 330294 158000 330914 187398
rect 334794 706758 335414 711590
rect 334794 706522 334826 706758
rect 335062 706522 335146 706758
rect 335382 706522 335414 706758
rect 334794 706438 335414 706522
rect 334794 706202 334826 706438
rect 335062 706202 335146 706438
rect 335382 706202 335414 706438
rect 334794 696454 335414 706202
rect 334794 696218 334826 696454
rect 335062 696218 335146 696454
rect 335382 696218 335414 696454
rect 334794 696134 335414 696218
rect 334794 695898 334826 696134
rect 335062 695898 335146 696134
rect 335382 695898 335414 696134
rect 334794 660454 335414 695898
rect 334794 660218 334826 660454
rect 335062 660218 335146 660454
rect 335382 660218 335414 660454
rect 334794 660134 335414 660218
rect 334794 659898 334826 660134
rect 335062 659898 335146 660134
rect 335382 659898 335414 660134
rect 334794 624454 335414 659898
rect 334794 624218 334826 624454
rect 335062 624218 335146 624454
rect 335382 624218 335414 624454
rect 334794 624134 335414 624218
rect 334794 623898 334826 624134
rect 335062 623898 335146 624134
rect 335382 623898 335414 624134
rect 334794 588454 335414 623898
rect 334794 588218 334826 588454
rect 335062 588218 335146 588454
rect 335382 588218 335414 588454
rect 334794 588134 335414 588218
rect 334794 587898 334826 588134
rect 335062 587898 335146 588134
rect 335382 587898 335414 588134
rect 334794 552454 335414 587898
rect 334794 552218 334826 552454
rect 335062 552218 335146 552454
rect 335382 552218 335414 552454
rect 334794 552134 335414 552218
rect 334794 551898 334826 552134
rect 335062 551898 335146 552134
rect 335382 551898 335414 552134
rect 334794 516454 335414 551898
rect 334794 516218 334826 516454
rect 335062 516218 335146 516454
rect 335382 516218 335414 516454
rect 334794 516134 335414 516218
rect 334794 515898 334826 516134
rect 335062 515898 335146 516134
rect 335382 515898 335414 516134
rect 334794 480454 335414 515898
rect 334794 480218 334826 480454
rect 335062 480218 335146 480454
rect 335382 480218 335414 480454
rect 334794 480134 335414 480218
rect 334794 479898 334826 480134
rect 335062 479898 335146 480134
rect 335382 479898 335414 480134
rect 334794 444454 335414 479898
rect 334794 444218 334826 444454
rect 335062 444218 335146 444454
rect 335382 444218 335414 444454
rect 334794 444134 335414 444218
rect 334794 443898 334826 444134
rect 335062 443898 335146 444134
rect 335382 443898 335414 444134
rect 334794 408454 335414 443898
rect 334794 408218 334826 408454
rect 335062 408218 335146 408454
rect 335382 408218 335414 408454
rect 334794 408134 335414 408218
rect 334794 407898 334826 408134
rect 335062 407898 335146 408134
rect 335382 407898 335414 408134
rect 334794 372454 335414 407898
rect 334794 372218 334826 372454
rect 335062 372218 335146 372454
rect 335382 372218 335414 372454
rect 334794 372134 335414 372218
rect 334794 371898 334826 372134
rect 335062 371898 335146 372134
rect 335382 371898 335414 372134
rect 334794 336454 335414 371898
rect 334794 336218 334826 336454
rect 335062 336218 335146 336454
rect 335382 336218 335414 336454
rect 334794 336134 335414 336218
rect 334794 335898 334826 336134
rect 335062 335898 335146 336134
rect 335382 335898 335414 336134
rect 334794 300454 335414 335898
rect 334794 300218 334826 300454
rect 335062 300218 335146 300454
rect 335382 300218 335414 300454
rect 334794 300134 335414 300218
rect 334794 299898 334826 300134
rect 335062 299898 335146 300134
rect 335382 299898 335414 300134
rect 334794 264454 335414 299898
rect 334794 264218 334826 264454
rect 335062 264218 335146 264454
rect 335382 264218 335414 264454
rect 334794 264134 335414 264218
rect 334794 263898 334826 264134
rect 335062 263898 335146 264134
rect 335382 263898 335414 264134
rect 334794 228454 335414 263898
rect 334794 228218 334826 228454
rect 335062 228218 335146 228454
rect 335382 228218 335414 228454
rect 334794 228134 335414 228218
rect 334794 227898 334826 228134
rect 335062 227898 335146 228134
rect 335382 227898 335414 228134
rect 334794 192454 335414 227898
rect 334794 192218 334826 192454
rect 335062 192218 335146 192454
rect 335382 192218 335414 192454
rect 334794 192134 335414 192218
rect 334794 191898 334826 192134
rect 335062 191898 335146 192134
rect 335382 191898 335414 192134
rect 334794 158000 335414 191898
rect 339294 707718 339914 711590
rect 339294 707482 339326 707718
rect 339562 707482 339646 707718
rect 339882 707482 339914 707718
rect 339294 707398 339914 707482
rect 339294 707162 339326 707398
rect 339562 707162 339646 707398
rect 339882 707162 339914 707398
rect 339294 700954 339914 707162
rect 339294 700718 339326 700954
rect 339562 700718 339646 700954
rect 339882 700718 339914 700954
rect 339294 700634 339914 700718
rect 339294 700398 339326 700634
rect 339562 700398 339646 700634
rect 339882 700398 339914 700634
rect 339294 664954 339914 700398
rect 339294 664718 339326 664954
rect 339562 664718 339646 664954
rect 339882 664718 339914 664954
rect 339294 664634 339914 664718
rect 339294 664398 339326 664634
rect 339562 664398 339646 664634
rect 339882 664398 339914 664634
rect 339294 628954 339914 664398
rect 339294 628718 339326 628954
rect 339562 628718 339646 628954
rect 339882 628718 339914 628954
rect 339294 628634 339914 628718
rect 339294 628398 339326 628634
rect 339562 628398 339646 628634
rect 339882 628398 339914 628634
rect 339294 592954 339914 628398
rect 339294 592718 339326 592954
rect 339562 592718 339646 592954
rect 339882 592718 339914 592954
rect 339294 592634 339914 592718
rect 339294 592398 339326 592634
rect 339562 592398 339646 592634
rect 339882 592398 339914 592634
rect 339294 556954 339914 592398
rect 339294 556718 339326 556954
rect 339562 556718 339646 556954
rect 339882 556718 339914 556954
rect 339294 556634 339914 556718
rect 339294 556398 339326 556634
rect 339562 556398 339646 556634
rect 339882 556398 339914 556634
rect 339294 520954 339914 556398
rect 339294 520718 339326 520954
rect 339562 520718 339646 520954
rect 339882 520718 339914 520954
rect 339294 520634 339914 520718
rect 339294 520398 339326 520634
rect 339562 520398 339646 520634
rect 339882 520398 339914 520634
rect 339294 484954 339914 520398
rect 339294 484718 339326 484954
rect 339562 484718 339646 484954
rect 339882 484718 339914 484954
rect 339294 484634 339914 484718
rect 339294 484398 339326 484634
rect 339562 484398 339646 484634
rect 339882 484398 339914 484634
rect 339294 448954 339914 484398
rect 339294 448718 339326 448954
rect 339562 448718 339646 448954
rect 339882 448718 339914 448954
rect 339294 448634 339914 448718
rect 339294 448398 339326 448634
rect 339562 448398 339646 448634
rect 339882 448398 339914 448634
rect 339294 412954 339914 448398
rect 339294 412718 339326 412954
rect 339562 412718 339646 412954
rect 339882 412718 339914 412954
rect 339294 412634 339914 412718
rect 339294 412398 339326 412634
rect 339562 412398 339646 412634
rect 339882 412398 339914 412634
rect 339294 376954 339914 412398
rect 343794 708678 344414 711590
rect 343794 708442 343826 708678
rect 344062 708442 344146 708678
rect 344382 708442 344414 708678
rect 343794 708358 344414 708442
rect 343794 708122 343826 708358
rect 344062 708122 344146 708358
rect 344382 708122 344414 708358
rect 343794 669454 344414 708122
rect 343794 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 344414 669454
rect 343794 669134 344414 669218
rect 343794 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 344414 669134
rect 343794 633454 344414 668898
rect 343794 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 344414 633454
rect 343794 633134 344414 633218
rect 343794 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 344414 633134
rect 343794 597454 344414 632898
rect 343794 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 344414 597454
rect 343794 597134 344414 597218
rect 343794 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 344414 597134
rect 343794 561454 344414 596898
rect 343794 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 344414 561454
rect 343794 561134 344414 561218
rect 343794 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 344414 561134
rect 343794 525454 344414 560898
rect 343794 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 344414 525454
rect 343794 525134 344414 525218
rect 343794 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 344414 525134
rect 343794 489454 344414 524898
rect 343794 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 344414 489454
rect 343794 489134 344414 489218
rect 343794 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 344414 489134
rect 343794 453454 344414 488898
rect 343794 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 344414 453454
rect 343794 453134 344414 453218
rect 343794 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 344414 453134
rect 343794 417454 344414 452898
rect 343794 417218 343826 417454
rect 344062 417218 344146 417454
rect 344382 417218 344414 417454
rect 343794 417134 344414 417218
rect 343794 416898 343826 417134
rect 344062 416898 344146 417134
rect 344382 416898 344414 417134
rect 342299 382804 342365 382805
rect 342299 382740 342300 382804
rect 342364 382740 342365 382804
rect 342299 382739 342365 382740
rect 339294 376718 339326 376954
rect 339562 376718 339646 376954
rect 339882 376718 339914 376954
rect 339294 376634 339914 376718
rect 339294 376398 339326 376634
rect 339562 376398 339646 376634
rect 339882 376398 339914 376634
rect 339294 340954 339914 376398
rect 339294 340718 339326 340954
rect 339562 340718 339646 340954
rect 339882 340718 339914 340954
rect 339294 340634 339914 340718
rect 339294 340398 339326 340634
rect 339562 340398 339646 340634
rect 339882 340398 339914 340634
rect 339294 304954 339914 340398
rect 339294 304718 339326 304954
rect 339562 304718 339646 304954
rect 339882 304718 339914 304954
rect 339294 304634 339914 304718
rect 339294 304398 339326 304634
rect 339562 304398 339646 304634
rect 339882 304398 339914 304634
rect 339294 268954 339914 304398
rect 339294 268718 339326 268954
rect 339562 268718 339646 268954
rect 339882 268718 339914 268954
rect 339294 268634 339914 268718
rect 339294 268398 339326 268634
rect 339562 268398 339646 268634
rect 339882 268398 339914 268634
rect 339294 232954 339914 268398
rect 339294 232718 339326 232954
rect 339562 232718 339646 232954
rect 339882 232718 339914 232954
rect 339294 232634 339914 232718
rect 339294 232398 339326 232634
rect 339562 232398 339646 232634
rect 339882 232398 339914 232634
rect 339294 196954 339914 232398
rect 339294 196718 339326 196954
rect 339562 196718 339646 196954
rect 339882 196718 339914 196954
rect 339294 196634 339914 196718
rect 339294 196398 339326 196634
rect 339562 196398 339646 196634
rect 339882 196398 339914 196634
rect 339294 160954 339914 196398
rect 339294 160718 339326 160954
rect 339562 160718 339646 160954
rect 339882 160718 339914 160954
rect 339294 160634 339914 160718
rect 339294 160398 339326 160634
rect 339562 160398 339646 160634
rect 339882 160398 339914 160634
rect 339294 158000 339914 160398
rect 284155 155684 284221 155685
rect 284155 155620 284156 155684
rect 284220 155620 284221 155684
rect 284155 155619 284221 155620
rect 296115 155684 296181 155685
rect 296115 155620 296116 155684
rect 296180 155620 296181 155684
rect 296115 155619 296181 155620
rect 270355 155548 270421 155549
rect 270355 155484 270356 155548
rect 270420 155484 270421 155548
rect 270355 155483 270421 155484
rect 284158 155277 284218 155619
rect 284155 155276 284221 155277
rect 284155 155212 284156 155276
rect 284220 155212 284221 155276
rect 284155 155211 284221 155212
rect 269067 153916 269133 153917
rect 269067 153852 269068 153916
rect 269132 153852 269133 153916
rect 269067 153851 269133 153852
rect 268147 153780 268213 153781
rect 268147 153716 268148 153780
rect 268212 153716 268213 153780
rect 268147 153715 268213 153716
rect 279568 151954 279888 151986
rect 279568 151718 279610 151954
rect 279846 151718 279888 151954
rect 279568 151634 279888 151718
rect 279568 151398 279610 151634
rect 279846 151398 279888 151634
rect 279568 151366 279888 151398
rect 310288 151954 310608 151986
rect 310288 151718 310330 151954
rect 310566 151718 310608 151954
rect 310288 151634 310608 151718
rect 310288 151398 310330 151634
rect 310566 151398 310608 151634
rect 310288 151366 310608 151398
rect 341008 151954 341328 151986
rect 341008 151718 341050 151954
rect 341286 151718 341328 151954
rect 341008 151634 341328 151718
rect 341008 151398 341050 151634
rect 341286 151398 341328 151634
rect 341008 151366 341328 151398
rect 264208 147454 264528 147486
rect 264208 147218 264250 147454
rect 264486 147218 264528 147454
rect 264208 147134 264528 147218
rect 264208 146898 264250 147134
rect 264486 146898 264528 147134
rect 264208 146866 264528 146898
rect 294928 147454 295248 147486
rect 294928 147218 294970 147454
rect 295206 147218 295248 147454
rect 294928 147134 295248 147218
rect 294928 146898 294970 147134
rect 295206 146898 295248 147134
rect 294928 146866 295248 146898
rect 325648 147454 325968 147486
rect 325648 147218 325690 147454
rect 325926 147218 325968 147454
rect 325648 147134 325968 147218
rect 325648 146898 325690 147134
rect 325926 146898 325968 147134
rect 325648 146866 325968 146898
rect 279568 115954 279888 115986
rect 279568 115718 279610 115954
rect 279846 115718 279888 115954
rect 279568 115634 279888 115718
rect 279568 115398 279610 115634
rect 279846 115398 279888 115634
rect 279568 115366 279888 115398
rect 310288 115954 310608 115986
rect 310288 115718 310330 115954
rect 310566 115718 310608 115954
rect 310288 115634 310608 115718
rect 310288 115398 310330 115634
rect 310566 115398 310608 115634
rect 310288 115366 310608 115398
rect 341008 115954 341328 115986
rect 341008 115718 341050 115954
rect 341286 115718 341328 115954
rect 341008 115634 341328 115718
rect 341008 115398 341050 115634
rect 341286 115398 341328 115634
rect 341008 115366 341328 115398
rect 264208 111454 264528 111486
rect 264208 111218 264250 111454
rect 264486 111218 264528 111454
rect 264208 111134 264528 111218
rect 264208 110898 264250 111134
rect 264486 110898 264528 111134
rect 264208 110866 264528 110898
rect 294928 111454 295248 111486
rect 294928 111218 294970 111454
rect 295206 111218 295248 111454
rect 294928 111134 295248 111218
rect 294928 110898 294970 111134
rect 295206 110898 295248 111134
rect 294928 110866 295248 110898
rect 325648 111454 325968 111486
rect 325648 111218 325690 111454
rect 325926 111218 325968 111454
rect 325648 111134 325968 111218
rect 325648 110898 325690 111134
rect 325926 110898 325968 111134
rect 325648 110866 325968 110898
rect 342302 100741 342362 382739
rect 342851 382668 342917 382669
rect 342851 382604 342852 382668
rect 342916 382604 342917 382668
rect 342851 382603 342917 382604
rect 342854 171150 342914 382603
rect 343794 381454 344414 416898
rect 348294 709638 348914 711590
rect 348294 709402 348326 709638
rect 348562 709402 348646 709638
rect 348882 709402 348914 709638
rect 348294 709318 348914 709402
rect 348294 709082 348326 709318
rect 348562 709082 348646 709318
rect 348882 709082 348914 709318
rect 348294 673954 348914 709082
rect 348294 673718 348326 673954
rect 348562 673718 348646 673954
rect 348882 673718 348914 673954
rect 348294 673634 348914 673718
rect 348294 673398 348326 673634
rect 348562 673398 348646 673634
rect 348882 673398 348914 673634
rect 348294 637954 348914 673398
rect 348294 637718 348326 637954
rect 348562 637718 348646 637954
rect 348882 637718 348914 637954
rect 348294 637634 348914 637718
rect 348294 637398 348326 637634
rect 348562 637398 348646 637634
rect 348882 637398 348914 637634
rect 348294 601954 348914 637398
rect 348294 601718 348326 601954
rect 348562 601718 348646 601954
rect 348882 601718 348914 601954
rect 348294 601634 348914 601718
rect 348294 601398 348326 601634
rect 348562 601398 348646 601634
rect 348882 601398 348914 601634
rect 348294 565954 348914 601398
rect 348294 565718 348326 565954
rect 348562 565718 348646 565954
rect 348882 565718 348914 565954
rect 348294 565634 348914 565718
rect 348294 565398 348326 565634
rect 348562 565398 348646 565634
rect 348882 565398 348914 565634
rect 348294 529954 348914 565398
rect 348294 529718 348326 529954
rect 348562 529718 348646 529954
rect 348882 529718 348914 529954
rect 348294 529634 348914 529718
rect 348294 529398 348326 529634
rect 348562 529398 348646 529634
rect 348882 529398 348914 529634
rect 348294 493954 348914 529398
rect 348294 493718 348326 493954
rect 348562 493718 348646 493954
rect 348882 493718 348914 493954
rect 348294 493634 348914 493718
rect 348294 493398 348326 493634
rect 348562 493398 348646 493634
rect 348882 493398 348914 493634
rect 348294 457954 348914 493398
rect 348294 457718 348326 457954
rect 348562 457718 348646 457954
rect 348882 457718 348914 457954
rect 348294 457634 348914 457718
rect 348294 457398 348326 457634
rect 348562 457398 348646 457634
rect 348882 457398 348914 457634
rect 348294 421954 348914 457398
rect 348294 421718 348326 421954
rect 348562 421718 348646 421954
rect 348882 421718 348914 421954
rect 348294 421634 348914 421718
rect 348294 421398 348326 421634
rect 348562 421398 348646 421634
rect 348882 421398 348914 421634
rect 348294 385954 348914 421398
rect 348294 385718 348326 385954
rect 348562 385718 348646 385954
rect 348882 385718 348914 385954
rect 348294 385634 348914 385718
rect 348294 385398 348326 385634
rect 348562 385398 348646 385634
rect 348882 385398 348914 385634
rect 345059 384300 345125 384301
rect 345059 384236 345060 384300
rect 345124 384236 345125 384300
rect 345059 384235 345125 384236
rect 343794 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 344414 381454
rect 343794 381134 344414 381218
rect 343794 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 344414 381134
rect 343794 345454 344414 380898
rect 343794 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 344414 345454
rect 343794 345134 344414 345218
rect 343794 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 344414 345134
rect 343794 309454 344414 344898
rect 344507 333844 344573 333845
rect 344507 333780 344508 333844
rect 344572 333780 344573 333844
rect 344507 333779 344573 333780
rect 343794 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 344414 309454
rect 343794 309134 344414 309218
rect 343794 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 344414 309134
rect 343794 273454 344414 308898
rect 343794 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 344414 273454
rect 343794 273134 344414 273218
rect 343794 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 344414 273134
rect 343794 237454 344414 272898
rect 343794 237218 343826 237454
rect 344062 237218 344146 237454
rect 344382 237218 344414 237454
rect 343794 237134 344414 237218
rect 343794 236898 343826 237134
rect 344062 236898 344146 237134
rect 344382 236898 344414 237134
rect 343794 201454 344414 236898
rect 343794 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 344414 201454
rect 343794 201134 344414 201218
rect 343794 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 344414 201134
rect 342854 171090 343466 171150
rect 343406 148341 343466 171090
rect 343794 165454 344414 200898
rect 343794 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 344414 165454
rect 343794 165134 344414 165218
rect 343794 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 344414 165134
rect 343587 161124 343653 161125
rect 343587 161060 343588 161124
rect 343652 161060 343653 161124
rect 343587 161059 343653 161060
rect 343403 148340 343469 148341
rect 343403 148276 343404 148340
rect 343468 148276 343469 148340
rect 343403 148275 343469 148276
rect 342299 100740 342365 100741
rect 342299 100676 342300 100740
rect 342364 100676 342365 100740
rect 342299 100675 342365 100676
rect 262794 84454 263414 98000
rect 262794 84218 262826 84454
rect 263062 84218 263146 84454
rect 263382 84218 263414 84454
rect 262794 84134 263414 84218
rect 262794 83898 262826 84134
rect 263062 83898 263146 84134
rect 263382 83898 263414 84134
rect 262794 48454 263414 83898
rect 262794 48218 262826 48454
rect 263062 48218 263146 48454
rect 263382 48218 263414 48454
rect 262794 48134 263414 48218
rect 262794 47898 262826 48134
rect 263062 47898 263146 48134
rect 263382 47898 263414 48134
rect 262794 12454 263414 47898
rect 262794 12218 262826 12454
rect 263062 12218 263146 12454
rect 263382 12218 263414 12454
rect 262794 12134 263414 12218
rect 262794 11898 262826 12134
rect 263062 11898 263146 12134
rect 263382 11898 263414 12134
rect 260603 3772 260669 3773
rect 260603 3708 260604 3772
rect 260668 3708 260669 3772
rect 260603 3707 260669 3708
rect 258294 -1542 258326 -1306
rect 258562 -1542 258646 -1306
rect 258882 -1542 258914 -1306
rect 258294 -1626 258914 -1542
rect 258294 -1862 258326 -1626
rect 258562 -1862 258646 -1626
rect 258882 -1862 258914 -1626
rect 258294 -7654 258914 -1862
rect 262794 -2266 263414 11898
rect 262794 -2502 262826 -2266
rect 263062 -2502 263146 -2266
rect 263382 -2502 263414 -2266
rect 262794 -2586 263414 -2502
rect 262794 -2822 262826 -2586
rect 263062 -2822 263146 -2586
rect 263382 -2822 263414 -2586
rect 262794 -7654 263414 -2822
rect 267294 88954 267914 98000
rect 267294 88718 267326 88954
rect 267562 88718 267646 88954
rect 267882 88718 267914 88954
rect 267294 88634 267914 88718
rect 267294 88398 267326 88634
rect 267562 88398 267646 88634
rect 267882 88398 267914 88634
rect 267294 52954 267914 88398
rect 267294 52718 267326 52954
rect 267562 52718 267646 52954
rect 267882 52718 267914 52954
rect 267294 52634 267914 52718
rect 267294 52398 267326 52634
rect 267562 52398 267646 52634
rect 267882 52398 267914 52634
rect 267294 16954 267914 52398
rect 267294 16718 267326 16954
rect 267562 16718 267646 16954
rect 267882 16718 267914 16954
rect 267294 16634 267914 16718
rect 267294 16398 267326 16634
rect 267562 16398 267646 16634
rect 267882 16398 267914 16634
rect 267294 -3226 267914 16398
rect 267294 -3462 267326 -3226
rect 267562 -3462 267646 -3226
rect 267882 -3462 267914 -3226
rect 267294 -3546 267914 -3462
rect 267294 -3782 267326 -3546
rect 267562 -3782 267646 -3546
rect 267882 -3782 267914 -3546
rect 267294 -7654 267914 -3782
rect 271794 93454 272414 98000
rect 271794 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 272414 93454
rect 271794 93134 272414 93218
rect 271794 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 272414 93134
rect 271794 57454 272414 92898
rect 271794 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 272414 57454
rect 271794 57134 272414 57218
rect 271794 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 272414 57134
rect 271794 21454 272414 56898
rect 271794 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 272414 21454
rect 271794 21134 272414 21218
rect 271794 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 272414 21134
rect 271794 -4186 272414 20898
rect 271794 -4422 271826 -4186
rect 272062 -4422 272146 -4186
rect 272382 -4422 272414 -4186
rect 271794 -4506 272414 -4422
rect 271794 -4742 271826 -4506
rect 272062 -4742 272146 -4506
rect 272382 -4742 272414 -4506
rect 271794 -7654 272414 -4742
rect 276294 97954 276914 98000
rect 276294 97718 276326 97954
rect 276562 97718 276646 97954
rect 276882 97718 276914 97954
rect 276294 97634 276914 97718
rect 276294 97398 276326 97634
rect 276562 97398 276646 97634
rect 276882 97398 276914 97634
rect 276294 61954 276914 97398
rect 276294 61718 276326 61954
rect 276562 61718 276646 61954
rect 276882 61718 276914 61954
rect 276294 61634 276914 61718
rect 276294 61398 276326 61634
rect 276562 61398 276646 61634
rect 276882 61398 276914 61634
rect 276294 25954 276914 61398
rect 276294 25718 276326 25954
rect 276562 25718 276646 25954
rect 276882 25718 276914 25954
rect 276294 25634 276914 25718
rect 276294 25398 276326 25634
rect 276562 25398 276646 25634
rect 276882 25398 276914 25634
rect 276294 -5146 276914 25398
rect 276294 -5382 276326 -5146
rect 276562 -5382 276646 -5146
rect 276882 -5382 276914 -5146
rect 276294 -5466 276914 -5382
rect 276294 -5702 276326 -5466
rect 276562 -5702 276646 -5466
rect 276882 -5702 276914 -5466
rect 276294 -7654 276914 -5702
rect 280794 66454 281414 98000
rect 280794 66218 280826 66454
rect 281062 66218 281146 66454
rect 281382 66218 281414 66454
rect 280794 66134 281414 66218
rect 280794 65898 280826 66134
rect 281062 65898 281146 66134
rect 281382 65898 281414 66134
rect 280794 30454 281414 65898
rect 280794 30218 280826 30454
rect 281062 30218 281146 30454
rect 281382 30218 281414 30454
rect 280794 30134 281414 30218
rect 280794 29898 280826 30134
rect 281062 29898 281146 30134
rect 281382 29898 281414 30134
rect 280794 -6106 281414 29898
rect 280794 -6342 280826 -6106
rect 281062 -6342 281146 -6106
rect 281382 -6342 281414 -6106
rect 280794 -6426 281414 -6342
rect 280794 -6662 280826 -6426
rect 281062 -6662 281146 -6426
rect 281382 -6662 281414 -6426
rect 280794 -7654 281414 -6662
rect 285294 70954 285914 98000
rect 285294 70718 285326 70954
rect 285562 70718 285646 70954
rect 285882 70718 285914 70954
rect 285294 70634 285914 70718
rect 285294 70398 285326 70634
rect 285562 70398 285646 70634
rect 285882 70398 285914 70634
rect 285294 34954 285914 70398
rect 285294 34718 285326 34954
rect 285562 34718 285646 34954
rect 285882 34718 285914 34954
rect 285294 34634 285914 34718
rect 285294 34398 285326 34634
rect 285562 34398 285646 34634
rect 285882 34398 285914 34634
rect 285294 -7066 285914 34398
rect 285294 -7302 285326 -7066
rect 285562 -7302 285646 -7066
rect 285882 -7302 285914 -7066
rect 285294 -7386 285914 -7302
rect 285294 -7622 285326 -7386
rect 285562 -7622 285646 -7386
rect 285882 -7622 285914 -7386
rect 285294 -7654 285914 -7622
rect 289794 75454 290414 98000
rect 289794 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 290414 75454
rect 289794 75134 290414 75218
rect 289794 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 290414 75134
rect 289794 39454 290414 74898
rect 289794 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 290414 39454
rect 289794 39134 290414 39218
rect 289794 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 290414 39134
rect 289794 3454 290414 38898
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -7654 290414 -902
rect 294294 79954 294914 98000
rect 294294 79718 294326 79954
rect 294562 79718 294646 79954
rect 294882 79718 294914 79954
rect 294294 79634 294914 79718
rect 294294 79398 294326 79634
rect 294562 79398 294646 79634
rect 294882 79398 294914 79634
rect 294294 43954 294914 79398
rect 294294 43718 294326 43954
rect 294562 43718 294646 43954
rect 294882 43718 294914 43954
rect 294294 43634 294914 43718
rect 294294 43398 294326 43634
rect 294562 43398 294646 43634
rect 294882 43398 294914 43634
rect 294294 7954 294914 43398
rect 294294 7718 294326 7954
rect 294562 7718 294646 7954
rect 294882 7718 294914 7954
rect 294294 7634 294914 7718
rect 294294 7398 294326 7634
rect 294562 7398 294646 7634
rect 294882 7398 294914 7634
rect 294294 -1306 294914 7398
rect 294294 -1542 294326 -1306
rect 294562 -1542 294646 -1306
rect 294882 -1542 294914 -1306
rect 294294 -1626 294914 -1542
rect 294294 -1862 294326 -1626
rect 294562 -1862 294646 -1626
rect 294882 -1862 294914 -1626
rect 294294 -7654 294914 -1862
rect 298794 84454 299414 98000
rect 298794 84218 298826 84454
rect 299062 84218 299146 84454
rect 299382 84218 299414 84454
rect 298794 84134 299414 84218
rect 298794 83898 298826 84134
rect 299062 83898 299146 84134
rect 299382 83898 299414 84134
rect 298794 48454 299414 83898
rect 298794 48218 298826 48454
rect 299062 48218 299146 48454
rect 299382 48218 299414 48454
rect 298794 48134 299414 48218
rect 298794 47898 298826 48134
rect 299062 47898 299146 48134
rect 299382 47898 299414 48134
rect 298794 12454 299414 47898
rect 298794 12218 298826 12454
rect 299062 12218 299146 12454
rect 299382 12218 299414 12454
rect 298794 12134 299414 12218
rect 298794 11898 298826 12134
rect 299062 11898 299146 12134
rect 299382 11898 299414 12134
rect 298794 -2266 299414 11898
rect 298794 -2502 298826 -2266
rect 299062 -2502 299146 -2266
rect 299382 -2502 299414 -2266
rect 298794 -2586 299414 -2502
rect 298794 -2822 298826 -2586
rect 299062 -2822 299146 -2586
rect 299382 -2822 299414 -2586
rect 298794 -7654 299414 -2822
rect 303294 88954 303914 98000
rect 303294 88718 303326 88954
rect 303562 88718 303646 88954
rect 303882 88718 303914 88954
rect 303294 88634 303914 88718
rect 303294 88398 303326 88634
rect 303562 88398 303646 88634
rect 303882 88398 303914 88634
rect 303294 52954 303914 88398
rect 303294 52718 303326 52954
rect 303562 52718 303646 52954
rect 303882 52718 303914 52954
rect 303294 52634 303914 52718
rect 303294 52398 303326 52634
rect 303562 52398 303646 52634
rect 303882 52398 303914 52634
rect 303294 16954 303914 52398
rect 303294 16718 303326 16954
rect 303562 16718 303646 16954
rect 303882 16718 303914 16954
rect 303294 16634 303914 16718
rect 303294 16398 303326 16634
rect 303562 16398 303646 16634
rect 303882 16398 303914 16634
rect 303294 -3226 303914 16398
rect 303294 -3462 303326 -3226
rect 303562 -3462 303646 -3226
rect 303882 -3462 303914 -3226
rect 303294 -3546 303914 -3462
rect 303294 -3782 303326 -3546
rect 303562 -3782 303646 -3546
rect 303882 -3782 303914 -3546
rect 303294 -7654 303914 -3782
rect 307794 93454 308414 98000
rect 307794 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 308414 93454
rect 307794 93134 308414 93218
rect 307794 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 308414 93134
rect 307794 57454 308414 92898
rect 307794 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 308414 57454
rect 307794 57134 308414 57218
rect 307794 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 308414 57134
rect 307794 21454 308414 56898
rect 307794 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 308414 21454
rect 307794 21134 308414 21218
rect 307794 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 308414 21134
rect 307794 -4186 308414 20898
rect 307794 -4422 307826 -4186
rect 308062 -4422 308146 -4186
rect 308382 -4422 308414 -4186
rect 307794 -4506 308414 -4422
rect 307794 -4742 307826 -4506
rect 308062 -4742 308146 -4506
rect 308382 -4742 308414 -4506
rect 307794 -7654 308414 -4742
rect 312294 97954 312914 98000
rect 312294 97718 312326 97954
rect 312562 97718 312646 97954
rect 312882 97718 312914 97954
rect 312294 97634 312914 97718
rect 312294 97398 312326 97634
rect 312562 97398 312646 97634
rect 312882 97398 312914 97634
rect 312294 61954 312914 97398
rect 312294 61718 312326 61954
rect 312562 61718 312646 61954
rect 312882 61718 312914 61954
rect 312294 61634 312914 61718
rect 312294 61398 312326 61634
rect 312562 61398 312646 61634
rect 312882 61398 312914 61634
rect 312294 25954 312914 61398
rect 312294 25718 312326 25954
rect 312562 25718 312646 25954
rect 312882 25718 312914 25954
rect 312294 25634 312914 25718
rect 312294 25398 312326 25634
rect 312562 25398 312646 25634
rect 312882 25398 312914 25634
rect 312294 -5146 312914 25398
rect 312294 -5382 312326 -5146
rect 312562 -5382 312646 -5146
rect 312882 -5382 312914 -5146
rect 312294 -5466 312914 -5382
rect 312294 -5702 312326 -5466
rect 312562 -5702 312646 -5466
rect 312882 -5702 312914 -5466
rect 312294 -7654 312914 -5702
rect 316794 66454 317414 98000
rect 316794 66218 316826 66454
rect 317062 66218 317146 66454
rect 317382 66218 317414 66454
rect 316794 66134 317414 66218
rect 316794 65898 316826 66134
rect 317062 65898 317146 66134
rect 317382 65898 317414 66134
rect 316794 30454 317414 65898
rect 316794 30218 316826 30454
rect 317062 30218 317146 30454
rect 317382 30218 317414 30454
rect 316794 30134 317414 30218
rect 316794 29898 316826 30134
rect 317062 29898 317146 30134
rect 317382 29898 317414 30134
rect 316794 -6106 317414 29898
rect 316794 -6342 316826 -6106
rect 317062 -6342 317146 -6106
rect 317382 -6342 317414 -6106
rect 316794 -6426 317414 -6342
rect 316794 -6662 316826 -6426
rect 317062 -6662 317146 -6426
rect 317382 -6662 317414 -6426
rect 316794 -7654 317414 -6662
rect 321294 70954 321914 98000
rect 321294 70718 321326 70954
rect 321562 70718 321646 70954
rect 321882 70718 321914 70954
rect 321294 70634 321914 70718
rect 321294 70398 321326 70634
rect 321562 70398 321646 70634
rect 321882 70398 321914 70634
rect 321294 34954 321914 70398
rect 321294 34718 321326 34954
rect 321562 34718 321646 34954
rect 321882 34718 321914 34954
rect 321294 34634 321914 34718
rect 321294 34398 321326 34634
rect 321562 34398 321646 34634
rect 321882 34398 321914 34634
rect 321294 -7066 321914 34398
rect 321294 -7302 321326 -7066
rect 321562 -7302 321646 -7066
rect 321882 -7302 321914 -7066
rect 321294 -7386 321914 -7302
rect 321294 -7622 321326 -7386
rect 321562 -7622 321646 -7386
rect 321882 -7622 321914 -7386
rect 321294 -7654 321914 -7622
rect 325794 75454 326414 98000
rect 325794 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 326414 75454
rect 325794 75134 326414 75218
rect 325794 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 326414 75134
rect 325794 39454 326414 74898
rect 325794 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 326414 39454
rect 325794 39134 326414 39218
rect 325794 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 326414 39134
rect 325794 3454 326414 38898
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -7654 326414 -902
rect 330294 79954 330914 98000
rect 330294 79718 330326 79954
rect 330562 79718 330646 79954
rect 330882 79718 330914 79954
rect 330294 79634 330914 79718
rect 330294 79398 330326 79634
rect 330562 79398 330646 79634
rect 330882 79398 330914 79634
rect 330294 43954 330914 79398
rect 330294 43718 330326 43954
rect 330562 43718 330646 43954
rect 330882 43718 330914 43954
rect 330294 43634 330914 43718
rect 330294 43398 330326 43634
rect 330562 43398 330646 43634
rect 330882 43398 330914 43634
rect 330294 7954 330914 43398
rect 330294 7718 330326 7954
rect 330562 7718 330646 7954
rect 330882 7718 330914 7954
rect 330294 7634 330914 7718
rect 330294 7398 330326 7634
rect 330562 7398 330646 7634
rect 330882 7398 330914 7634
rect 330294 -1306 330914 7398
rect 330294 -1542 330326 -1306
rect 330562 -1542 330646 -1306
rect 330882 -1542 330914 -1306
rect 330294 -1626 330914 -1542
rect 330294 -1862 330326 -1626
rect 330562 -1862 330646 -1626
rect 330882 -1862 330914 -1626
rect 330294 -7654 330914 -1862
rect 334794 84454 335414 98000
rect 334794 84218 334826 84454
rect 335062 84218 335146 84454
rect 335382 84218 335414 84454
rect 334794 84134 335414 84218
rect 334794 83898 334826 84134
rect 335062 83898 335146 84134
rect 335382 83898 335414 84134
rect 334794 48454 335414 83898
rect 334794 48218 334826 48454
rect 335062 48218 335146 48454
rect 335382 48218 335414 48454
rect 334794 48134 335414 48218
rect 334794 47898 334826 48134
rect 335062 47898 335146 48134
rect 335382 47898 335414 48134
rect 334794 12454 335414 47898
rect 334794 12218 334826 12454
rect 335062 12218 335146 12454
rect 335382 12218 335414 12454
rect 334794 12134 335414 12218
rect 334794 11898 334826 12134
rect 335062 11898 335146 12134
rect 335382 11898 335414 12134
rect 334794 -2266 335414 11898
rect 334794 -2502 334826 -2266
rect 335062 -2502 335146 -2266
rect 335382 -2502 335414 -2266
rect 334794 -2586 335414 -2502
rect 334794 -2822 334826 -2586
rect 335062 -2822 335146 -2586
rect 335382 -2822 335414 -2586
rect 334794 -7654 335414 -2822
rect 339294 88954 339914 98000
rect 339294 88718 339326 88954
rect 339562 88718 339646 88954
rect 339882 88718 339914 88954
rect 339294 88634 339914 88718
rect 339294 88398 339326 88634
rect 339562 88398 339646 88634
rect 339882 88398 339914 88634
rect 339294 52954 339914 88398
rect 339294 52718 339326 52954
rect 339562 52718 339646 52954
rect 339882 52718 339914 52954
rect 339294 52634 339914 52718
rect 339294 52398 339326 52634
rect 339562 52398 339646 52634
rect 339882 52398 339914 52634
rect 339294 16954 339914 52398
rect 339294 16718 339326 16954
rect 339562 16718 339646 16954
rect 339882 16718 339914 16954
rect 339294 16634 339914 16718
rect 339294 16398 339326 16634
rect 339562 16398 339646 16634
rect 339882 16398 339914 16634
rect 339294 -3226 339914 16398
rect 343590 3501 343650 161059
rect 343794 158000 344414 164898
rect 343794 93454 344414 98000
rect 343794 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 344414 93454
rect 343794 93134 344414 93218
rect 343794 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 344414 93134
rect 343794 57454 344414 92898
rect 343794 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 344414 57454
rect 343794 57134 344414 57218
rect 343794 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 344414 57134
rect 343794 21454 344414 56898
rect 343794 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 344414 21454
rect 343794 21134 344414 21218
rect 343794 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 344414 21134
rect 343587 3500 343653 3501
rect 343587 3436 343588 3500
rect 343652 3436 343653 3500
rect 343587 3435 343653 3436
rect 339294 -3462 339326 -3226
rect 339562 -3462 339646 -3226
rect 339882 -3462 339914 -3226
rect 339294 -3546 339914 -3462
rect 339294 -3782 339326 -3546
rect 339562 -3782 339646 -3546
rect 339882 -3782 339914 -3546
rect 339294 -7654 339914 -3782
rect 343794 -4186 344414 20898
rect 344510 3090 344570 333779
rect 344691 157452 344757 157453
rect 344691 157388 344692 157452
rect 344756 157388 344757 157452
rect 344691 157387 344757 157388
rect 344694 129845 344754 157387
rect 344691 129844 344757 129845
rect 344691 129780 344692 129844
rect 344756 129780 344757 129844
rect 344691 129779 344757 129780
rect 345062 97885 345122 384235
rect 345243 381852 345309 381853
rect 345243 381788 345244 381852
rect 345308 381788 345309 381852
rect 345243 381787 345309 381788
rect 345246 142901 345306 381787
rect 346899 381444 346965 381445
rect 346899 381380 346900 381444
rect 346964 381380 346965 381444
rect 346899 381379 346965 381380
rect 345427 161396 345493 161397
rect 345427 161332 345428 161396
rect 345492 161332 345493 161396
rect 345427 161331 345493 161332
rect 345243 142900 345309 142901
rect 345243 142836 345244 142900
rect 345308 142836 345309 142900
rect 345243 142835 345309 142836
rect 345430 121141 345490 161331
rect 345427 121140 345493 121141
rect 345427 121076 345428 121140
rect 345492 121076 345493 121140
rect 345427 121075 345493 121076
rect 345059 97884 345125 97885
rect 345059 97820 345060 97884
rect 345124 97820 345125 97884
rect 345059 97819 345125 97820
rect 346902 31789 346962 381379
rect 348294 349954 348914 385398
rect 348294 349718 348326 349954
rect 348562 349718 348646 349954
rect 348882 349718 348914 349954
rect 348294 349634 348914 349718
rect 348294 349398 348326 349634
rect 348562 349398 348646 349634
rect 348882 349398 348914 349634
rect 348294 313954 348914 349398
rect 348294 313718 348326 313954
rect 348562 313718 348646 313954
rect 348882 313718 348914 313954
rect 348294 313634 348914 313718
rect 348294 313398 348326 313634
rect 348562 313398 348646 313634
rect 348882 313398 348914 313634
rect 348294 277954 348914 313398
rect 348294 277718 348326 277954
rect 348562 277718 348646 277954
rect 348882 277718 348914 277954
rect 348294 277634 348914 277718
rect 348294 277398 348326 277634
rect 348562 277398 348646 277634
rect 348882 277398 348914 277634
rect 348294 241954 348914 277398
rect 348294 241718 348326 241954
rect 348562 241718 348646 241954
rect 348882 241718 348914 241954
rect 348294 241634 348914 241718
rect 348294 241398 348326 241634
rect 348562 241398 348646 241634
rect 348882 241398 348914 241634
rect 348294 205954 348914 241398
rect 348294 205718 348326 205954
rect 348562 205718 348646 205954
rect 348882 205718 348914 205954
rect 348294 205634 348914 205718
rect 348294 205398 348326 205634
rect 348562 205398 348646 205634
rect 348882 205398 348914 205634
rect 348294 169954 348914 205398
rect 348294 169718 348326 169954
rect 348562 169718 348646 169954
rect 348882 169718 348914 169954
rect 348294 169634 348914 169718
rect 348294 169398 348326 169634
rect 348562 169398 348646 169634
rect 348882 169398 348914 169634
rect 348294 133954 348914 169398
rect 348294 133718 348326 133954
rect 348562 133718 348646 133954
rect 348882 133718 348914 133954
rect 348294 133634 348914 133718
rect 348294 133398 348326 133634
rect 348562 133398 348646 133634
rect 348882 133398 348914 133634
rect 348294 97954 348914 133398
rect 348294 97718 348326 97954
rect 348562 97718 348646 97954
rect 348882 97718 348914 97954
rect 348294 97634 348914 97718
rect 348294 97398 348326 97634
rect 348562 97398 348646 97634
rect 348882 97398 348914 97634
rect 348294 61954 348914 97398
rect 348294 61718 348326 61954
rect 348562 61718 348646 61954
rect 348882 61718 348914 61954
rect 348294 61634 348914 61718
rect 348294 61398 348326 61634
rect 348562 61398 348646 61634
rect 348882 61398 348914 61634
rect 346899 31788 346965 31789
rect 346899 31724 346900 31788
rect 346964 31724 346965 31788
rect 346899 31723 346965 31724
rect 348294 25954 348914 61398
rect 348294 25718 348326 25954
rect 348562 25718 348646 25954
rect 348882 25718 348914 25954
rect 348294 25634 348914 25718
rect 348294 25398 348326 25634
rect 348562 25398 348646 25634
rect 348882 25398 348914 25634
rect 344967 3228 345033 3229
rect 344967 3164 344968 3228
rect 345032 3164 345033 3228
rect 344967 3163 345033 3164
rect 344970 3090 345030 3163
rect 344510 3030 345030 3090
rect 343794 -4422 343826 -4186
rect 344062 -4422 344146 -4186
rect 344382 -4422 344414 -4186
rect 343794 -4506 344414 -4422
rect 343794 -4742 343826 -4506
rect 344062 -4742 344146 -4506
rect 344382 -4742 344414 -4506
rect 343794 -7654 344414 -4742
rect 348294 -5146 348914 25398
rect 348294 -5382 348326 -5146
rect 348562 -5382 348646 -5146
rect 348882 -5382 348914 -5146
rect 348294 -5466 348914 -5382
rect 348294 -5702 348326 -5466
rect 348562 -5702 348646 -5466
rect 348882 -5702 348914 -5466
rect 348294 -7654 348914 -5702
rect 352794 710598 353414 711590
rect 352794 710362 352826 710598
rect 353062 710362 353146 710598
rect 353382 710362 353414 710598
rect 352794 710278 353414 710362
rect 352794 710042 352826 710278
rect 353062 710042 353146 710278
rect 353382 710042 353414 710278
rect 352794 678454 353414 710042
rect 352794 678218 352826 678454
rect 353062 678218 353146 678454
rect 353382 678218 353414 678454
rect 352794 678134 353414 678218
rect 352794 677898 352826 678134
rect 353062 677898 353146 678134
rect 353382 677898 353414 678134
rect 352794 642454 353414 677898
rect 352794 642218 352826 642454
rect 353062 642218 353146 642454
rect 353382 642218 353414 642454
rect 352794 642134 353414 642218
rect 352794 641898 352826 642134
rect 353062 641898 353146 642134
rect 353382 641898 353414 642134
rect 352794 606454 353414 641898
rect 352794 606218 352826 606454
rect 353062 606218 353146 606454
rect 353382 606218 353414 606454
rect 352794 606134 353414 606218
rect 352794 605898 352826 606134
rect 353062 605898 353146 606134
rect 353382 605898 353414 606134
rect 352794 570454 353414 605898
rect 352794 570218 352826 570454
rect 353062 570218 353146 570454
rect 353382 570218 353414 570454
rect 352794 570134 353414 570218
rect 352794 569898 352826 570134
rect 353062 569898 353146 570134
rect 353382 569898 353414 570134
rect 352794 534454 353414 569898
rect 352794 534218 352826 534454
rect 353062 534218 353146 534454
rect 353382 534218 353414 534454
rect 352794 534134 353414 534218
rect 352794 533898 352826 534134
rect 353062 533898 353146 534134
rect 353382 533898 353414 534134
rect 352794 498454 353414 533898
rect 352794 498218 352826 498454
rect 353062 498218 353146 498454
rect 353382 498218 353414 498454
rect 352794 498134 353414 498218
rect 352794 497898 352826 498134
rect 353062 497898 353146 498134
rect 353382 497898 353414 498134
rect 352794 462454 353414 497898
rect 352794 462218 352826 462454
rect 353062 462218 353146 462454
rect 353382 462218 353414 462454
rect 352794 462134 353414 462218
rect 352794 461898 352826 462134
rect 353062 461898 353146 462134
rect 353382 461898 353414 462134
rect 352794 426454 353414 461898
rect 352794 426218 352826 426454
rect 353062 426218 353146 426454
rect 353382 426218 353414 426454
rect 352794 426134 353414 426218
rect 352794 425898 352826 426134
rect 353062 425898 353146 426134
rect 353382 425898 353414 426134
rect 352794 390454 353414 425898
rect 352794 390218 352826 390454
rect 353062 390218 353146 390454
rect 353382 390218 353414 390454
rect 352794 390134 353414 390218
rect 352794 389898 352826 390134
rect 353062 389898 353146 390134
rect 353382 389898 353414 390134
rect 352794 354454 353414 389898
rect 352794 354218 352826 354454
rect 353062 354218 353146 354454
rect 353382 354218 353414 354454
rect 352794 354134 353414 354218
rect 352794 353898 352826 354134
rect 353062 353898 353146 354134
rect 353382 353898 353414 354134
rect 352794 318454 353414 353898
rect 352794 318218 352826 318454
rect 353062 318218 353146 318454
rect 353382 318218 353414 318454
rect 352794 318134 353414 318218
rect 352794 317898 352826 318134
rect 353062 317898 353146 318134
rect 353382 317898 353414 318134
rect 352794 282454 353414 317898
rect 352794 282218 352826 282454
rect 353062 282218 353146 282454
rect 353382 282218 353414 282454
rect 352794 282134 353414 282218
rect 352794 281898 352826 282134
rect 353062 281898 353146 282134
rect 353382 281898 353414 282134
rect 352794 246454 353414 281898
rect 352794 246218 352826 246454
rect 353062 246218 353146 246454
rect 353382 246218 353414 246454
rect 352794 246134 353414 246218
rect 352794 245898 352826 246134
rect 353062 245898 353146 246134
rect 353382 245898 353414 246134
rect 352794 210454 353414 245898
rect 352794 210218 352826 210454
rect 353062 210218 353146 210454
rect 353382 210218 353414 210454
rect 352794 210134 353414 210218
rect 352794 209898 352826 210134
rect 353062 209898 353146 210134
rect 353382 209898 353414 210134
rect 352794 174454 353414 209898
rect 352794 174218 352826 174454
rect 353062 174218 353146 174454
rect 353382 174218 353414 174454
rect 352794 174134 353414 174218
rect 352794 173898 352826 174134
rect 353062 173898 353146 174134
rect 353382 173898 353414 174134
rect 352794 138454 353414 173898
rect 352794 138218 352826 138454
rect 353062 138218 353146 138454
rect 353382 138218 353414 138454
rect 352794 138134 353414 138218
rect 352794 137898 352826 138134
rect 353062 137898 353146 138134
rect 353382 137898 353414 138134
rect 352794 102454 353414 137898
rect 352794 102218 352826 102454
rect 353062 102218 353146 102454
rect 353382 102218 353414 102454
rect 352794 102134 353414 102218
rect 352794 101898 352826 102134
rect 353062 101898 353146 102134
rect 353382 101898 353414 102134
rect 352794 66454 353414 101898
rect 352794 66218 352826 66454
rect 353062 66218 353146 66454
rect 353382 66218 353414 66454
rect 352794 66134 353414 66218
rect 352794 65898 352826 66134
rect 353062 65898 353146 66134
rect 353382 65898 353414 66134
rect 352794 30454 353414 65898
rect 352794 30218 352826 30454
rect 353062 30218 353146 30454
rect 353382 30218 353414 30454
rect 352794 30134 353414 30218
rect 352794 29898 352826 30134
rect 353062 29898 353146 30134
rect 353382 29898 353414 30134
rect 352794 -6106 353414 29898
rect 352794 -6342 352826 -6106
rect 353062 -6342 353146 -6106
rect 353382 -6342 353414 -6106
rect 352794 -6426 353414 -6342
rect 352794 -6662 352826 -6426
rect 353062 -6662 353146 -6426
rect 353382 -6662 353414 -6426
rect 352794 -7654 353414 -6662
rect 357294 711558 357914 711590
rect 357294 711322 357326 711558
rect 357562 711322 357646 711558
rect 357882 711322 357914 711558
rect 357294 711238 357914 711322
rect 357294 711002 357326 711238
rect 357562 711002 357646 711238
rect 357882 711002 357914 711238
rect 357294 682954 357914 711002
rect 357294 682718 357326 682954
rect 357562 682718 357646 682954
rect 357882 682718 357914 682954
rect 357294 682634 357914 682718
rect 357294 682398 357326 682634
rect 357562 682398 357646 682634
rect 357882 682398 357914 682634
rect 357294 646954 357914 682398
rect 357294 646718 357326 646954
rect 357562 646718 357646 646954
rect 357882 646718 357914 646954
rect 357294 646634 357914 646718
rect 357294 646398 357326 646634
rect 357562 646398 357646 646634
rect 357882 646398 357914 646634
rect 357294 610954 357914 646398
rect 357294 610718 357326 610954
rect 357562 610718 357646 610954
rect 357882 610718 357914 610954
rect 357294 610634 357914 610718
rect 357294 610398 357326 610634
rect 357562 610398 357646 610634
rect 357882 610398 357914 610634
rect 357294 574954 357914 610398
rect 357294 574718 357326 574954
rect 357562 574718 357646 574954
rect 357882 574718 357914 574954
rect 357294 574634 357914 574718
rect 357294 574398 357326 574634
rect 357562 574398 357646 574634
rect 357882 574398 357914 574634
rect 357294 538954 357914 574398
rect 357294 538718 357326 538954
rect 357562 538718 357646 538954
rect 357882 538718 357914 538954
rect 357294 538634 357914 538718
rect 357294 538398 357326 538634
rect 357562 538398 357646 538634
rect 357882 538398 357914 538634
rect 357294 502954 357914 538398
rect 357294 502718 357326 502954
rect 357562 502718 357646 502954
rect 357882 502718 357914 502954
rect 357294 502634 357914 502718
rect 357294 502398 357326 502634
rect 357562 502398 357646 502634
rect 357882 502398 357914 502634
rect 357294 466954 357914 502398
rect 357294 466718 357326 466954
rect 357562 466718 357646 466954
rect 357882 466718 357914 466954
rect 357294 466634 357914 466718
rect 357294 466398 357326 466634
rect 357562 466398 357646 466634
rect 357882 466398 357914 466634
rect 357294 430954 357914 466398
rect 357294 430718 357326 430954
rect 357562 430718 357646 430954
rect 357882 430718 357914 430954
rect 357294 430634 357914 430718
rect 357294 430398 357326 430634
rect 357562 430398 357646 430634
rect 357882 430398 357914 430634
rect 357294 394954 357914 430398
rect 357294 394718 357326 394954
rect 357562 394718 357646 394954
rect 357882 394718 357914 394954
rect 357294 394634 357914 394718
rect 357294 394398 357326 394634
rect 357562 394398 357646 394634
rect 357882 394398 357914 394634
rect 357294 358954 357914 394398
rect 357294 358718 357326 358954
rect 357562 358718 357646 358954
rect 357882 358718 357914 358954
rect 357294 358634 357914 358718
rect 357294 358398 357326 358634
rect 357562 358398 357646 358634
rect 357882 358398 357914 358634
rect 357294 322954 357914 358398
rect 357294 322718 357326 322954
rect 357562 322718 357646 322954
rect 357882 322718 357914 322954
rect 357294 322634 357914 322718
rect 357294 322398 357326 322634
rect 357562 322398 357646 322634
rect 357882 322398 357914 322634
rect 357294 286954 357914 322398
rect 357294 286718 357326 286954
rect 357562 286718 357646 286954
rect 357882 286718 357914 286954
rect 357294 286634 357914 286718
rect 357294 286398 357326 286634
rect 357562 286398 357646 286634
rect 357882 286398 357914 286634
rect 357294 250954 357914 286398
rect 357294 250718 357326 250954
rect 357562 250718 357646 250954
rect 357882 250718 357914 250954
rect 357294 250634 357914 250718
rect 357294 250398 357326 250634
rect 357562 250398 357646 250634
rect 357882 250398 357914 250634
rect 357294 214954 357914 250398
rect 357294 214718 357326 214954
rect 357562 214718 357646 214954
rect 357882 214718 357914 214954
rect 357294 214634 357914 214718
rect 357294 214398 357326 214634
rect 357562 214398 357646 214634
rect 357882 214398 357914 214634
rect 357294 178954 357914 214398
rect 357294 178718 357326 178954
rect 357562 178718 357646 178954
rect 357882 178718 357914 178954
rect 357294 178634 357914 178718
rect 357294 178398 357326 178634
rect 357562 178398 357646 178634
rect 357882 178398 357914 178634
rect 357294 142954 357914 178398
rect 357294 142718 357326 142954
rect 357562 142718 357646 142954
rect 357882 142718 357914 142954
rect 357294 142634 357914 142718
rect 357294 142398 357326 142634
rect 357562 142398 357646 142634
rect 357882 142398 357914 142634
rect 357294 106954 357914 142398
rect 357294 106718 357326 106954
rect 357562 106718 357646 106954
rect 357882 106718 357914 106954
rect 357294 106634 357914 106718
rect 357294 106398 357326 106634
rect 357562 106398 357646 106634
rect 357882 106398 357914 106634
rect 357294 70954 357914 106398
rect 357294 70718 357326 70954
rect 357562 70718 357646 70954
rect 357882 70718 357914 70954
rect 357294 70634 357914 70718
rect 357294 70398 357326 70634
rect 357562 70398 357646 70634
rect 357882 70398 357914 70634
rect 357294 34954 357914 70398
rect 357294 34718 357326 34954
rect 357562 34718 357646 34954
rect 357882 34718 357914 34954
rect 357294 34634 357914 34718
rect 357294 34398 357326 34634
rect 357562 34398 357646 34634
rect 357882 34398 357914 34634
rect 357294 -7066 357914 34398
rect 357294 -7302 357326 -7066
rect 357562 -7302 357646 -7066
rect 357882 -7302 357914 -7066
rect 357294 -7386 357914 -7302
rect 357294 -7622 357326 -7386
rect 357562 -7622 357646 -7386
rect 357882 -7622 357914 -7386
rect 357294 -7654 357914 -7622
rect 361794 704838 362414 711590
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 687454 362414 704282
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 361794 651454 362414 686898
rect 361794 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 362414 651454
rect 361794 651134 362414 651218
rect 361794 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 362414 651134
rect 361794 615454 362414 650898
rect 361794 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 362414 615454
rect 361794 615134 362414 615218
rect 361794 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 362414 615134
rect 361794 579454 362414 614898
rect 361794 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 362414 579454
rect 361794 579134 362414 579218
rect 361794 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 362414 579134
rect 361794 543454 362414 578898
rect 361794 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 362414 543454
rect 361794 543134 362414 543218
rect 361794 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 362414 543134
rect 361794 507454 362414 542898
rect 361794 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 362414 507454
rect 361794 507134 362414 507218
rect 361794 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 362414 507134
rect 361794 471454 362414 506898
rect 361794 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 362414 471454
rect 361794 471134 362414 471218
rect 361794 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 362414 471134
rect 361794 435454 362414 470898
rect 361794 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 362414 435454
rect 361794 435134 362414 435218
rect 361794 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 362414 435134
rect 361794 399454 362414 434898
rect 361794 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 362414 399454
rect 361794 399134 362414 399218
rect 361794 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 362414 399134
rect 361794 363454 362414 398898
rect 361794 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 362414 363454
rect 361794 363134 362414 363218
rect 361794 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 362414 363134
rect 361794 327454 362414 362898
rect 361794 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 362414 327454
rect 361794 327134 362414 327218
rect 361794 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 362414 327134
rect 361794 291454 362414 326898
rect 361794 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 362414 291454
rect 361794 291134 362414 291218
rect 361794 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 362414 291134
rect 361794 255454 362414 290898
rect 361794 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 362414 255454
rect 361794 255134 362414 255218
rect 361794 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 362414 255134
rect 361794 219454 362414 254898
rect 361794 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 362414 219454
rect 361794 219134 362414 219218
rect 361794 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 362414 219134
rect 361794 183454 362414 218898
rect 361794 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 362414 183454
rect 361794 183134 362414 183218
rect 361794 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 362414 183134
rect 361794 147454 362414 182898
rect 361794 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 362414 147454
rect 361794 147134 362414 147218
rect 361794 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 362414 147134
rect 361794 111454 362414 146898
rect 361794 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 362414 111454
rect 361794 111134 362414 111218
rect 361794 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 362414 111134
rect 361794 75454 362414 110898
rect 361794 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 362414 75454
rect 361794 75134 362414 75218
rect 361794 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 362414 75134
rect 361794 39454 362414 74898
rect 361794 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 362414 39454
rect 361794 39134 362414 39218
rect 361794 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 362414 39134
rect 361794 3454 362414 38898
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -7654 362414 -902
rect 366294 705798 366914 711590
rect 366294 705562 366326 705798
rect 366562 705562 366646 705798
rect 366882 705562 366914 705798
rect 366294 705478 366914 705562
rect 366294 705242 366326 705478
rect 366562 705242 366646 705478
rect 366882 705242 366914 705478
rect 366294 691954 366914 705242
rect 366294 691718 366326 691954
rect 366562 691718 366646 691954
rect 366882 691718 366914 691954
rect 366294 691634 366914 691718
rect 366294 691398 366326 691634
rect 366562 691398 366646 691634
rect 366882 691398 366914 691634
rect 366294 655954 366914 691398
rect 366294 655718 366326 655954
rect 366562 655718 366646 655954
rect 366882 655718 366914 655954
rect 366294 655634 366914 655718
rect 366294 655398 366326 655634
rect 366562 655398 366646 655634
rect 366882 655398 366914 655634
rect 366294 619954 366914 655398
rect 366294 619718 366326 619954
rect 366562 619718 366646 619954
rect 366882 619718 366914 619954
rect 366294 619634 366914 619718
rect 366294 619398 366326 619634
rect 366562 619398 366646 619634
rect 366882 619398 366914 619634
rect 366294 583954 366914 619398
rect 366294 583718 366326 583954
rect 366562 583718 366646 583954
rect 366882 583718 366914 583954
rect 366294 583634 366914 583718
rect 366294 583398 366326 583634
rect 366562 583398 366646 583634
rect 366882 583398 366914 583634
rect 366294 547954 366914 583398
rect 366294 547718 366326 547954
rect 366562 547718 366646 547954
rect 366882 547718 366914 547954
rect 366294 547634 366914 547718
rect 366294 547398 366326 547634
rect 366562 547398 366646 547634
rect 366882 547398 366914 547634
rect 366294 511954 366914 547398
rect 366294 511718 366326 511954
rect 366562 511718 366646 511954
rect 366882 511718 366914 511954
rect 366294 511634 366914 511718
rect 366294 511398 366326 511634
rect 366562 511398 366646 511634
rect 366882 511398 366914 511634
rect 366294 475954 366914 511398
rect 366294 475718 366326 475954
rect 366562 475718 366646 475954
rect 366882 475718 366914 475954
rect 366294 475634 366914 475718
rect 366294 475398 366326 475634
rect 366562 475398 366646 475634
rect 366882 475398 366914 475634
rect 366294 439954 366914 475398
rect 366294 439718 366326 439954
rect 366562 439718 366646 439954
rect 366882 439718 366914 439954
rect 366294 439634 366914 439718
rect 366294 439398 366326 439634
rect 366562 439398 366646 439634
rect 366882 439398 366914 439634
rect 366294 403954 366914 439398
rect 366294 403718 366326 403954
rect 366562 403718 366646 403954
rect 366882 403718 366914 403954
rect 366294 403634 366914 403718
rect 366294 403398 366326 403634
rect 366562 403398 366646 403634
rect 366882 403398 366914 403634
rect 366294 367954 366914 403398
rect 366294 367718 366326 367954
rect 366562 367718 366646 367954
rect 366882 367718 366914 367954
rect 366294 367634 366914 367718
rect 366294 367398 366326 367634
rect 366562 367398 366646 367634
rect 366882 367398 366914 367634
rect 366294 331954 366914 367398
rect 366294 331718 366326 331954
rect 366562 331718 366646 331954
rect 366882 331718 366914 331954
rect 366294 331634 366914 331718
rect 366294 331398 366326 331634
rect 366562 331398 366646 331634
rect 366882 331398 366914 331634
rect 366294 295954 366914 331398
rect 366294 295718 366326 295954
rect 366562 295718 366646 295954
rect 366882 295718 366914 295954
rect 366294 295634 366914 295718
rect 366294 295398 366326 295634
rect 366562 295398 366646 295634
rect 366882 295398 366914 295634
rect 366294 259954 366914 295398
rect 366294 259718 366326 259954
rect 366562 259718 366646 259954
rect 366882 259718 366914 259954
rect 366294 259634 366914 259718
rect 366294 259398 366326 259634
rect 366562 259398 366646 259634
rect 366882 259398 366914 259634
rect 366294 223954 366914 259398
rect 366294 223718 366326 223954
rect 366562 223718 366646 223954
rect 366882 223718 366914 223954
rect 366294 223634 366914 223718
rect 366294 223398 366326 223634
rect 366562 223398 366646 223634
rect 366882 223398 366914 223634
rect 366294 187954 366914 223398
rect 366294 187718 366326 187954
rect 366562 187718 366646 187954
rect 366882 187718 366914 187954
rect 366294 187634 366914 187718
rect 366294 187398 366326 187634
rect 366562 187398 366646 187634
rect 366882 187398 366914 187634
rect 366294 151954 366914 187398
rect 366294 151718 366326 151954
rect 366562 151718 366646 151954
rect 366882 151718 366914 151954
rect 366294 151634 366914 151718
rect 366294 151398 366326 151634
rect 366562 151398 366646 151634
rect 366882 151398 366914 151634
rect 366294 115954 366914 151398
rect 366294 115718 366326 115954
rect 366562 115718 366646 115954
rect 366882 115718 366914 115954
rect 366294 115634 366914 115718
rect 366294 115398 366326 115634
rect 366562 115398 366646 115634
rect 366882 115398 366914 115634
rect 366294 79954 366914 115398
rect 366294 79718 366326 79954
rect 366562 79718 366646 79954
rect 366882 79718 366914 79954
rect 366294 79634 366914 79718
rect 366294 79398 366326 79634
rect 366562 79398 366646 79634
rect 366882 79398 366914 79634
rect 366294 43954 366914 79398
rect 366294 43718 366326 43954
rect 366562 43718 366646 43954
rect 366882 43718 366914 43954
rect 366294 43634 366914 43718
rect 366294 43398 366326 43634
rect 366562 43398 366646 43634
rect 366882 43398 366914 43634
rect 366294 7954 366914 43398
rect 366294 7718 366326 7954
rect 366562 7718 366646 7954
rect 366882 7718 366914 7954
rect 366294 7634 366914 7718
rect 366294 7398 366326 7634
rect 366562 7398 366646 7634
rect 366882 7398 366914 7634
rect 366294 -1306 366914 7398
rect 366294 -1542 366326 -1306
rect 366562 -1542 366646 -1306
rect 366882 -1542 366914 -1306
rect 366294 -1626 366914 -1542
rect 366294 -1862 366326 -1626
rect 366562 -1862 366646 -1626
rect 366882 -1862 366914 -1626
rect 366294 -7654 366914 -1862
rect 370794 706758 371414 711590
rect 370794 706522 370826 706758
rect 371062 706522 371146 706758
rect 371382 706522 371414 706758
rect 370794 706438 371414 706522
rect 370794 706202 370826 706438
rect 371062 706202 371146 706438
rect 371382 706202 371414 706438
rect 370794 696454 371414 706202
rect 370794 696218 370826 696454
rect 371062 696218 371146 696454
rect 371382 696218 371414 696454
rect 370794 696134 371414 696218
rect 370794 695898 370826 696134
rect 371062 695898 371146 696134
rect 371382 695898 371414 696134
rect 370794 660454 371414 695898
rect 370794 660218 370826 660454
rect 371062 660218 371146 660454
rect 371382 660218 371414 660454
rect 370794 660134 371414 660218
rect 370794 659898 370826 660134
rect 371062 659898 371146 660134
rect 371382 659898 371414 660134
rect 370794 624454 371414 659898
rect 370794 624218 370826 624454
rect 371062 624218 371146 624454
rect 371382 624218 371414 624454
rect 370794 624134 371414 624218
rect 370794 623898 370826 624134
rect 371062 623898 371146 624134
rect 371382 623898 371414 624134
rect 370794 588454 371414 623898
rect 370794 588218 370826 588454
rect 371062 588218 371146 588454
rect 371382 588218 371414 588454
rect 370794 588134 371414 588218
rect 370794 587898 370826 588134
rect 371062 587898 371146 588134
rect 371382 587898 371414 588134
rect 370794 552454 371414 587898
rect 370794 552218 370826 552454
rect 371062 552218 371146 552454
rect 371382 552218 371414 552454
rect 370794 552134 371414 552218
rect 370794 551898 370826 552134
rect 371062 551898 371146 552134
rect 371382 551898 371414 552134
rect 370794 516454 371414 551898
rect 370794 516218 370826 516454
rect 371062 516218 371146 516454
rect 371382 516218 371414 516454
rect 370794 516134 371414 516218
rect 370794 515898 370826 516134
rect 371062 515898 371146 516134
rect 371382 515898 371414 516134
rect 370794 480454 371414 515898
rect 370794 480218 370826 480454
rect 371062 480218 371146 480454
rect 371382 480218 371414 480454
rect 370794 480134 371414 480218
rect 370794 479898 370826 480134
rect 371062 479898 371146 480134
rect 371382 479898 371414 480134
rect 370794 444454 371414 479898
rect 370794 444218 370826 444454
rect 371062 444218 371146 444454
rect 371382 444218 371414 444454
rect 370794 444134 371414 444218
rect 370794 443898 370826 444134
rect 371062 443898 371146 444134
rect 371382 443898 371414 444134
rect 370794 408454 371414 443898
rect 370794 408218 370826 408454
rect 371062 408218 371146 408454
rect 371382 408218 371414 408454
rect 370794 408134 371414 408218
rect 370794 407898 370826 408134
rect 371062 407898 371146 408134
rect 371382 407898 371414 408134
rect 370794 372454 371414 407898
rect 370794 372218 370826 372454
rect 371062 372218 371146 372454
rect 371382 372218 371414 372454
rect 370794 372134 371414 372218
rect 370794 371898 370826 372134
rect 371062 371898 371146 372134
rect 371382 371898 371414 372134
rect 370794 336454 371414 371898
rect 370794 336218 370826 336454
rect 371062 336218 371146 336454
rect 371382 336218 371414 336454
rect 370794 336134 371414 336218
rect 370794 335898 370826 336134
rect 371062 335898 371146 336134
rect 371382 335898 371414 336134
rect 370794 300454 371414 335898
rect 370794 300218 370826 300454
rect 371062 300218 371146 300454
rect 371382 300218 371414 300454
rect 370794 300134 371414 300218
rect 370794 299898 370826 300134
rect 371062 299898 371146 300134
rect 371382 299898 371414 300134
rect 370794 264454 371414 299898
rect 370794 264218 370826 264454
rect 371062 264218 371146 264454
rect 371382 264218 371414 264454
rect 370794 264134 371414 264218
rect 370794 263898 370826 264134
rect 371062 263898 371146 264134
rect 371382 263898 371414 264134
rect 370794 228454 371414 263898
rect 370794 228218 370826 228454
rect 371062 228218 371146 228454
rect 371382 228218 371414 228454
rect 370794 228134 371414 228218
rect 370794 227898 370826 228134
rect 371062 227898 371146 228134
rect 371382 227898 371414 228134
rect 370794 192454 371414 227898
rect 370794 192218 370826 192454
rect 371062 192218 371146 192454
rect 371382 192218 371414 192454
rect 370794 192134 371414 192218
rect 370794 191898 370826 192134
rect 371062 191898 371146 192134
rect 371382 191898 371414 192134
rect 370794 156454 371414 191898
rect 370794 156218 370826 156454
rect 371062 156218 371146 156454
rect 371382 156218 371414 156454
rect 370794 156134 371414 156218
rect 370794 155898 370826 156134
rect 371062 155898 371146 156134
rect 371382 155898 371414 156134
rect 370794 120454 371414 155898
rect 370794 120218 370826 120454
rect 371062 120218 371146 120454
rect 371382 120218 371414 120454
rect 370794 120134 371414 120218
rect 370794 119898 370826 120134
rect 371062 119898 371146 120134
rect 371382 119898 371414 120134
rect 370794 84454 371414 119898
rect 370794 84218 370826 84454
rect 371062 84218 371146 84454
rect 371382 84218 371414 84454
rect 370794 84134 371414 84218
rect 370794 83898 370826 84134
rect 371062 83898 371146 84134
rect 371382 83898 371414 84134
rect 370794 48454 371414 83898
rect 370794 48218 370826 48454
rect 371062 48218 371146 48454
rect 371382 48218 371414 48454
rect 370794 48134 371414 48218
rect 370794 47898 370826 48134
rect 371062 47898 371146 48134
rect 371382 47898 371414 48134
rect 370794 12454 371414 47898
rect 370794 12218 370826 12454
rect 371062 12218 371146 12454
rect 371382 12218 371414 12454
rect 370794 12134 371414 12218
rect 370794 11898 370826 12134
rect 371062 11898 371146 12134
rect 371382 11898 371414 12134
rect 370794 -2266 371414 11898
rect 370794 -2502 370826 -2266
rect 371062 -2502 371146 -2266
rect 371382 -2502 371414 -2266
rect 370794 -2586 371414 -2502
rect 370794 -2822 370826 -2586
rect 371062 -2822 371146 -2586
rect 371382 -2822 371414 -2586
rect 370794 -7654 371414 -2822
rect 375294 707718 375914 711590
rect 375294 707482 375326 707718
rect 375562 707482 375646 707718
rect 375882 707482 375914 707718
rect 375294 707398 375914 707482
rect 375294 707162 375326 707398
rect 375562 707162 375646 707398
rect 375882 707162 375914 707398
rect 375294 700954 375914 707162
rect 375294 700718 375326 700954
rect 375562 700718 375646 700954
rect 375882 700718 375914 700954
rect 375294 700634 375914 700718
rect 375294 700398 375326 700634
rect 375562 700398 375646 700634
rect 375882 700398 375914 700634
rect 375294 664954 375914 700398
rect 375294 664718 375326 664954
rect 375562 664718 375646 664954
rect 375882 664718 375914 664954
rect 375294 664634 375914 664718
rect 375294 664398 375326 664634
rect 375562 664398 375646 664634
rect 375882 664398 375914 664634
rect 375294 628954 375914 664398
rect 375294 628718 375326 628954
rect 375562 628718 375646 628954
rect 375882 628718 375914 628954
rect 375294 628634 375914 628718
rect 375294 628398 375326 628634
rect 375562 628398 375646 628634
rect 375882 628398 375914 628634
rect 375294 592954 375914 628398
rect 375294 592718 375326 592954
rect 375562 592718 375646 592954
rect 375882 592718 375914 592954
rect 375294 592634 375914 592718
rect 375294 592398 375326 592634
rect 375562 592398 375646 592634
rect 375882 592398 375914 592634
rect 375294 556954 375914 592398
rect 379794 708678 380414 711590
rect 379794 708442 379826 708678
rect 380062 708442 380146 708678
rect 380382 708442 380414 708678
rect 379794 708358 380414 708442
rect 379794 708122 379826 708358
rect 380062 708122 380146 708358
rect 380382 708122 380414 708358
rect 379794 669454 380414 708122
rect 379794 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 380414 669454
rect 379794 669134 380414 669218
rect 379794 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 380414 669134
rect 379794 633454 380414 668898
rect 379794 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 380414 633454
rect 379794 633134 380414 633218
rect 379794 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 380414 633134
rect 379794 597454 380414 632898
rect 379794 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 380414 597454
rect 379794 597134 380414 597218
rect 379794 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 380414 597134
rect 379794 591292 380414 596898
rect 384294 709638 384914 711590
rect 384294 709402 384326 709638
rect 384562 709402 384646 709638
rect 384882 709402 384914 709638
rect 384294 709318 384914 709402
rect 384294 709082 384326 709318
rect 384562 709082 384646 709318
rect 384882 709082 384914 709318
rect 384294 673954 384914 709082
rect 384294 673718 384326 673954
rect 384562 673718 384646 673954
rect 384882 673718 384914 673954
rect 384294 673634 384914 673718
rect 384294 673398 384326 673634
rect 384562 673398 384646 673634
rect 384882 673398 384914 673634
rect 384294 637954 384914 673398
rect 384294 637718 384326 637954
rect 384562 637718 384646 637954
rect 384882 637718 384914 637954
rect 384294 637634 384914 637718
rect 384294 637398 384326 637634
rect 384562 637398 384646 637634
rect 384882 637398 384914 637634
rect 384294 601954 384914 637398
rect 384294 601718 384326 601954
rect 384562 601718 384646 601954
rect 384882 601718 384914 601954
rect 384294 601634 384914 601718
rect 384294 601398 384326 601634
rect 384562 601398 384646 601634
rect 384882 601398 384914 601634
rect 384294 591292 384914 601398
rect 388794 710598 389414 711590
rect 388794 710362 388826 710598
rect 389062 710362 389146 710598
rect 389382 710362 389414 710598
rect 388794 710278 389414 710362
rect 388794 710042 388826 710278
rect 389062 710042 389146 710278
rect 389382 710042 389414 710278
rect 388794 678454 389414 710042
rect 388794 678218 388826 678454
rect 389062 678218 389146 678454
rect 389382 678218 389414 678454
rect 388794 678134 389414 678218
rect 388794 677898 388826 678134
rect 389062 677898 389146 678134
rect 389382 677898 389414 678134
rect 388794 642454 389414 677898
rect 388794 642218 388826 642454
rect 389062 642218 389146 642454
rect 389382 642218 389414 642454
rect 388794 642134 389414 642218
rect 388794 641898 388826 642134
rect 389062 641898 389146 642134
rect 389382 641898 389414 642134
rect 388794 606454 389414 641898
rect 388794 606218 388826 606454
rect 389062 606218 389146 606454
rect 389382 606218 389414 606454
rect 388794 606134 389414 606218
rect 388794 605898 388826 606134
rect 389062 605898 389146 606134
rect 389382 605898 389414 606134
rect 388794 591292 389414 605898
rect 393294 711558 393914 711590
rect 393294 711322 393326 711558
rect 393562 711322 393646 711558
rect 393882 711322 393914 711558
rect 393294 711238 393914 711322
rect 393294 711002 393326 711238
rect 393562 711002 393646 711238
rect 393882 711002 393914 711238
rect 393294 682954 393914 711002
rect 393294 682718 393326 682954
rect 393562 682718 393646 682954
rect 393882 682718 393914 682954
rect 393294 682634 393914 682718
rect 393294 682398 393326 682634
rect 393562 682398 393646 682634
rect 393882 682398 393914 682634
rect 393294 646954 393914 682398
rect 393294 646718 393326 646954
rect 393562 646718 393646 646954
rect 393882 646718 393914 646954
rect 393294 646634 393914 646718
rect 393294 646398 393326 646634
rect 393562 646398 393646 646634
rect 393882 646398 393914 646634
rect 393294 610954 393914 646398
rect 393294 610718 393326 610954
rect 393562 610718 393646 610954
rect 393882 610718 393914 610954
rect 393294 610634 393914 610718
rect 393294 610398 393326 610634
rect 393562 610398 393646 610634
rect 393882 610398 393914 610634
rect 393294 591292 393914 610398
rect 397794 704838 398414 711590
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 687454 398414 704282
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 651454 398414 686898
rect 397794 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 398414 651454
rect 397794 651134 398414 651218
rect 397794 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 398414 651134
rect 397794 615454 398414 650898
rect 397794 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 398414 615454
rect 397794 615134 398414 615218
rect 397794 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 398414 615134
rect 397794 591292 398414 614898
rect 402294 705798 402914 711590
rect 402294 705562 402326 705798
rect 402562 705562 402646 705798
rect 402882 705562 402914 705798
rect 402294 705478 402914 705562
rect 402294 705242 402326 705478
rect 402562 705242 402646 705478
rect 402882 705242 402914 705478
rect 402294 691954 402914 705242
rect 402294 691718 402326 691954
rect 402562 691718 402646 691954
rect 402882 691718 402914 691954
rect 402294 691634 402914 691718
rect 402294 691398 402326 691634
rect 402562 691398 402646 691634
rect 402882 691398 402914 691634
rect 402294 655954 402914 691398
rect 402294 655718 402326 655954
rect 402562 655718 402646 655954
rect 402882 655718 402914 655954
rect 402294 655634 402914 655718
rect 402294 655398 402326 655634
rect 402562 655398 402646 655634
rect 402882 655398 402914 655634
rect 402294 619954 402914 655398
rect 402294 619718 402326 619954
rect 402562 619718 402646 619954
rect 402882 619718 402914 619954
rect 402294 619634 402914 619718
rect 402294 619398 402326 619634
rect 402562 619398 402646 619634
rect 402882 619398 402914 619634
rect 402294 591292 402914 619398
rect 406794 706758 407414 711590
rect 406794 706522 406826 706758
rect 407062 706522 407146 706758
rect 407382 706522 407414 706758
rect 406794 706438 407414 706522
rect 406794 706202 406826 706438
rect 407062 706202 407146 706438
rect 407382 706202 407414 706438
rect 406794 696454 407414 706202
rect 406794 696218 406826 696454
rect 407062 696218 407146 696454
rect 407382 696218 407414 696454
rect 406794 696134 407414 696218
rect 406794 695898 406826 696134
rect 407062 695898 407146 696134
rect 407382 695898 407414 696134
rect 406794 660454 407414 695898
rect 406794 660218 406826 660454
rect 407062 660218 407146 660454
rect 407382 660218 407414 660454
rect 406794 660134 407414 660218
rect 406794 659898 406826 660134
rect 407062 659898 407146 660134
rect 407382 659898 407414 660134
rect 406794 624454 407414 659898
rect 406794 624218 406826 624454
rect 407062 624218 407146 624454
rect 407382 624218 407414 624454
rect 406794 624134 407414 624218
rect 406794 623898 406826 624134
rect 407062 623898 407146 624134
rect 407382 623898 407414 624134
rect 406794 591292 407414 623898
rect 411294 707718 411914 711590
rect 411294 707482 411326 707718
rect 411562 707482 411646 707718
rect 411882 707482 411914 707718
rect 411294 707398 411914 707482
rect 411294 707162 411326 707398
rect 411562 707162 411646 707398
rect 411882 707162 411914 707398
rect 411294 700954 411914 707162
rect 411294 700718 411326 700954
rect 411562 700718 411646 700954
rect 411882 700718 411914 700954
rect 411294 700634 411914 700718
rect 411294 700398 411326 700634
rect 411562 700398 411646 700634
rect 411882 700398 411914 700634
rect 411294 664954 411914 700398
rect 411294 664718 411326 664954
rect 411562 664718 411646 664954
rect 411882 664718 411914 664954
rect 411294 664634 411914 664718
rect 411294 664398 411326 664634
rect 411562 664398 411646 664634
rect 411882 664398 411914 664634
rect 411294 628954 411914 664398
rect 411294 628718 411326 628954
rect 411562 628718 411646 628954
rect 411882 628718 411914 628954
rect 411294 628634 411914 628718
rect 411294 628398 411326 628634
rect 411562 628398 411646 628634
rect 411882 628398 411914 628634
rect 411294 592954 411914 628398
rect 411294 592718 411326 592954
rect 411562 592718 411646 592954
rect 411882 592718 411914 592954
rect 411294 592634 411914 592718
rect 411294 592398 411326 592634
rect 411562 592398 411646 592634
rect 411882 592398 411914 592634
rect 411294 591292 411914 592398
rect 415794 708678 416414 711590
rect 415794 708442 415826 708678
rect 416062 708442 416146 708678
rect 416382 708442 416414 708678
rect 415794 708358 416414 708442
rect 415794 708122 415826 708358
rect 416062 708122 416146 708358
rect 416382 708122 416414 708358
rect 415794 669454 416414 708122
rect 415794 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 416414 669454
rect 415794 669134 416414 669218
rect 415794 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 416414 669134
rect 415794 633454 416414 668898
rect 415794 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 416414 633454
rect 415794 633134 416414 633218
rect 415794 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 416414 633134
rect 415794 597454 416414 632898
rect 415794 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 416414 597454
rect 415794 597134 416414 597218
rect 415794 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 416414 597134
rect 415794 591292 416414 596898
rect 420294 709638 420914 711590
rect 420294 709402 420326 709638
rect 420562 709402 420646 709638
rect 420882 709402 420914 709638
rect 420294 709318 420914 709402
rect 420294 709082 420326 709318
rect 420562 709082 420646 709318
rect 420882 709082 420914 709318
rect 420294 673954 420914 709082
rect 420294 673718 420326 673954
rect 420562 673718 420646 673954
rect 420882 673718 420914 673954
rect 420294 673634 420914 673718
rect 420294 673398 420326 673634
rect 420562 673398 420646 673634
rect 420882 673398 420914 673634
rect 420294 637954 420914 673398
rect 420294 637718 420326 637954
rect 420562 637718 420646 637954
rect 420882 637718 420914 637954
rect 420294 637634 420914 637718
rect 420294 637398 420326 637634
rect 420562 637398 420646 637634
rect 420882 637398 420914 637634
rect 420294 601954 420914 637398
rect 420294 601718 420326 601954
rect 420562 601718 420646 601954
rect 420882 601718 420914 601954
rect 420294 601634 420914 601718
rect 420294 601398 420326 601634
rect 420562 601398 420646 601634
rect 420882 601398 420914 601634
rect 420294 591292 420914 601398
rect 424794 710598 425414 711590
rect 424794 710362 424826 710598
rect 425062 710362 425146 710598
rect 425382 710362 425414 710598
rect 424794 710278 425414 710362
rect 424794 710042 424826 710278
rect 425062 710042 425146 710278
rect 425382 710042 425414 710278
rect 424794 678454 425414 710042
rect 424794 678218 424826 678454
rect 425062 678218 425146 678454
rect 425382 678218 425414 678454
rect 424794 678134 425414 678218
rect 424794 677898 424826 678134
rect 425062 677898 425146 678134
rect 425382 677898 425414 678134
rect 424794 642454 425414 677898
rect 424794 642218 424826 642454
rect 425062 642218 425146 642454
rect 425382 642218 425414 642454
rect 424794 642134 425414 642218
rect 424794 641898 424826 642134
rect 425062 641898 425146 642134
rect 425382 641898 425414 642134
rect 424794 606454 425414 641898
rect 424794 606218 424826 606454
rect 425062 606218 425146 606454
rect 425382 606218 425414 606454
rect 424794 606134 425414 606218
rect 424794 605898 424826 606134
rect 425062 605898 425146 606134
rect 425382 605898 425414 606134
rect 424794 591292 425414 605898
rect 429294 711558 429914 711590
rect 429294 711322 429326 711558
rect 429562 711322 429646 711558
rect 429882 711322 429914 711558
rect 429294 711238 429914 711322
rect 429294 711002 429326 711238
rect 429562 711002 429646 711238
rect 429882 711002 429914 711238
rect 429294 682954 429914 711002
rect 429294 682718 429326 682954
rect 429562 682718 429646 682954
rect 429882 682718 429914 682954
rect 429294 682634 429914 682718
rect 429294 682398 429326 682634
rect 429562 682398 429646 682634
rect 429882 682398 429914 682634
rect 429294 646954 429914 682398
rect 429294 646718 429326 646954
rect 429562 646718 429646 646954
rect 429882 646718 429914 646954
rect 429294 646634 429914 646718
rect 429294 646398 429326 646634
rect 429562 646398 429646 646634
rect 429882 646398 429914 646634
rect 429294 610954 429914 646398
rect 429294 610718 429326 610954
rect 429562 610718 429646 610954
rect 429882 610718 429914 610954
rect 429294 610634 429914 610718
rect 429294 610398 429326 610634
rect 429562 610398 429646 610634
rect 429882 610398 429914 610634
rect 429294 591292 429914 610398
rect 433794 704838 434414 711590
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 687454 434414 704282
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 651454 434414 686898
rect 433794 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 434414 651454
rect 433794 651134 434414 651218
rect 433794 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 434414 651134
rect 433794 615454 434414 650898
rect 433794 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 434414 615454
rect 433794 615134 434414 615218
rect 433794 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 434414 615134
rect 433794 591292 434414 614898
rect 438294 705798 438914 711590
rect 438294 705562 438326 705798
rect 438562 705562 438646 705798
rect 438882 705562 438914 705798
rect 438294 705478 438914 705562
rect 438294 705242 438326 705478
rect 438562 705242 438646 705478
rect 438882 705242 438914 705478
rect 438294 691954 438914 705242
rect 438294 691718 438326 691954
rect 438562 691718 438646 691954
rect 438882 691718 438914 691954
rect 438294 691634 438914 691718
rect 438294 691398 438326 691634
rect 438562 691398 438646 691634
rect 438882 691398 438914 691634
rect 438294 655954 438914 691398
rect 438294 655718 438326 655954
rect 438562 655718 438646 655954
rect 438882 655718 438914 655954
rect 438294 655634 438914 655718
rect 438294 655398 438326 655634
rect 438562 655398 438646 655634
rect 438882 655398 438914 655634
rect 438294 619954 438914 655398
rect 438294 619718 438326 619954
rect 438562 619718 438646 619954
rect 438882 619718 438914 619954
rect 438294 619634 438914 619718
rect 438294 619398 438326 619634
rect 438562 619398 438646 619634
rect 438882 619398 438914 619634
rect 438294 591292 438914 619398
rect 442794 706758 443414 711590
rect 442794 706522 442826 706758
rect 443062 706522 443146 706758
rect 443382 706522 443414 706758
rect 442794 706438 443414 706522
rect 442794 706202 442826 706438
rect 443062 706202 443146 706438
rect 443382 706202 443414 706438
rect 442794 696454 443414 706202
rect 442794 696218 442826 696454
rect 443062 696218 443146 696454
rect 443382 696218 443414 696454
rect 442794 696134 443414 696218
rect 442794 695898 442826 696134
rect 443062 695898 443146 696134
rect 443382 695898 443414 696134
rect 442794 660454 443414 695898
rect 442794 660218 442826 660454
rect 443062 660218 443146 660454
rect 443382 660218 443414 660454
rect 442794 660134 443414 660218
rect 442794 659898 442826 660134
rect 443062 659898 443146 660134
rect 443382 659898 443414 660134
rect 442794 624454 443414 659898
rect 442794 624218 442826 624454
rect 443062 624218 443146 624454
rect 443382 624218 443414 624454
rect 442794 624134 443414 624218
rect 442794 623898 442826 624134
rect 443062 623898 443146 624134
rect 443382 623898 443414 624134
rect 442794 591292 443414 623898
rect 447294 707718 447914 711590
rect 447294 707482 447326 707718
rect 447562 707482 447646 707718
rect 447882 707482 447914 707718
rect 447294 707398 447914 707482
rect 447294 707162 447326 707398
rect 447562 707162 447646 707398
rect 447882 707162 447914 707398
rect 447294 700954 447914 707162
rect 447294 700718 447326 700954
rect 447562 700718 447646 700954
rect 447882 700718 447914 700954
rect 447294 700634 447914 700718
rect 447294 700398 447326 700634
rect 447562 700398 447646 700634
rect 447882 700398 447914 700634
rect 447294 664954 447914 700398
rect 447294 664718 447326 664954
rect 447562 664718 447646 664954
rect 447882 664718 447914 664954
rect 447294 664634 447914 664718
rect 447294 664398 447326 664634
rect 447562 664398 447646 664634
rect 447882 664398 447914 664634
rect 447294 628954 447914 664398
rect 447294 628718 447326 628954
rect 447562 628718 447646 628954
rect 447882 628718 447914 628954
rect 447294 628634 447914 628718
rect 447294 628398 447326 628634
rect 447562 628398 447646 628634
rect 447882 628398 447914 628634
rect 447294 592954 447914 628398
rect 447294 592718 447326 592954
rect 447562 592718 447646 592954
rect 447882 592718 447914 592954
rect 447294 592634 447914 592718
rect 447294 592398 447326 592634
rect 447562 592398 447646 592634
rect 447882 592398 447914 592634
rect 447294 591292 447914 592398
rect 451794 708678 452414 711590
rect 451794 708442 451826 708678
rect 452062 708442 452146 708678
rect 452382 708442 452414 708678
rect 451794 708358 452414 708442
rect 451794 708122 451826 708358
rect 452062 708122 452146 708358
rect 452382 708122 452414 708358
rect 451794 669454 452414 708122
rect 451794 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 452414 669454
rect 451794 669134 452414 669218
rect 451794 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 452414 669134
rect 451794 633454 452414 668898
rect 451794 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 452414 633454
rect 451794 633134 452414 633218
rect 451794 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 452414 633134
rect 451794 597454 452414 632898
rect 451794 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 452414 597454
rect 451794 597134 452414 597218
rect 451794 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 452414 597134
rect 451794 591292 452414 596898
rect 456294 709638 456914 711590
rect 456294 709402 456326 709638
rect 456562 709402 456646 709638
rect 456882 709402 456914 709638
rect 456294 709318 456914 709402
rect 456294 709082 456326 709318
rect 456562 709082 456646 709318
rect 456882 709082 456914 709318
rect 456294 673954 456914 709082
rect 456294 673718 456326 673954
rect 456562 673718 456646 673954
rect 456882 673718 456914 673954
rect 456294 673634 456914 673718
rect 456294 673398 456326 673634
rect 456562 673398 456646 673634
rect 456882 673398 456914 673634
rect 456294 637954 456914 673398
rect 456294 637718 456326 637954
rect 456562 637718 456646 637954
rect 456882 637718 456914 637954
rect 456294 637634 456914 637718
rect 456294 637398 456326 637634
rect 456562 637398 456646 637634
rect 456882 637398 456914 637634
rect 456294 601954 456914 637398
rect 456294 601718 456326 601954
rect 456562 601718 456646 601954
rect 456882 601718 456914 601954
rect 456294 601634 456914 601718
rect 456294 601398 456326 601634
rect 456562 601398 456646 601634
rect 456882 601398 456914 601634
rect 456294 591292 456914 601398
rect 460794 710598 461414 711590
rect 460794 710362 460826 710598
rect 461062 710362 461146 710598
rect 461382 710362 461414 710598
rect 460794 710278 461414 710362
rect 460794 710042 460826 710278
rect 461062 710042 461146 710278
rect 461382 710042 461414 710278
rect 460794 678454 461414 710042
rect 460794 678218 460826 678454
rect 461062 678218 461146 678454
rect 461382 678218 461414 678454
rect 460794 678134 461414 678218
rect 460794 677898 460826 678134
rect 461062 677898 461146 678134
rect 461382 677898 461414 678134
rect 460794 642454 461414 677898
rect 460794 642218 460826 642454
rect 461062 642218 461146 642454
rect 461382 642218 461414 642454
rect 460794 642134 461414 642218
rect 460794 641898 460826 642134
rect 461062 641898 461146 642134
rect 461382 641898 461414 642134
rect 460794 606454 461414 641898
rect 460794 606218 460826 606454
rect 461062 606218 461146 606454
rect 461382 606218 461414 606454
rect 460794 606134 461414 606218
rect 460794 605898 460826 606134
rect 461062 605898 461146 606134
rect 461382 605898 461414 606134
rect 460794 591292 461414 605898
rect 465294 711558 465914 711590
rect 465294 711322 465326 711558
rect 465562 711322 465646 711558
rect 465882 711322 465914 711558
rect 465294 711238 465914 711322
rect 465294 711002 465326 711238
rect 465562 711002 465646 711238
rect 465882 711002 465914 711238
rect 465294 682954 465914 711002
rect 465294 682718 465326 682954
rect 465562 682718 465646 682954
rect 465882 682718 465914 682954
rect 465294 682634 465914 682718
rect 465294 682398 465326 682634
rect 465562 682398 465646 682634
rect 465882 682398 465914 682634
rect 465294 646954 465914 682398
rect 465294 646718 465326 646954
rect 465562 646718 465646 646954
rect 465882 646718 465914 646954
rect 465294 646634 465914 646718
rect 465294 646398 465326 646634
rect 465562 646398 465646 646634
rect 465882 646398 465914 646634
rect 465294 610954 465914 646398
rect 465294 610718 465326 610954
rect 465562 610718 465646 610954
rect 465882 610718 465914 610954
rect 465294 610634 465914 610718
rect 465294 610398 465326 610634
rect 465562 610398 465646 610634
rect 465882 610398 465914 610634
rect 465294 591292 465914 610398
rect 469794 704838 470414 711590
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 687454 470414 704282
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469794 651454 470414 686898
rect 469794 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 470414 651454
rect 469794 651134 470414 651218
rect 469794 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 470414 651134
rect 469794 615454 470414 650898
rect 469794 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 470414 615454
rect 469794 615134 470414 615218
rect 469794 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 470414 615134
rect 469794 591292 470414 614898
rect 474294 705798 474914 711590
rect 474294 705562 474326 705798
rect 474562 705562 474646 705798
rect 474882 705562 474914 705798
rect 474294 705478 474914 705562
rect 474294 705242 474326 705478
rect 474562 705242 474646 705478
rect 474882 705242 474914 705478
rect 474294 691954 474914 705242
rect 474294 691718 474326 691954
rect 474562 691718 474646 691954
rect 474882 691718 474914 691954
rect 474294 691634 474914 691718
rect 474294 691398 474326 691634
rect 474562 691398 474646 691634
rect 474882 691398 474914 691634
rect 474294 655954 474914 691398
rect 474294 655718 474326 655954
rect 474562 655718 474646 655954
rect 474882 655718 474914 655954
rect 474294 655634 474914 655718
rect 474294 655398 474326 655634
rect 474562 655398 474646 655634
rect 474882 655398 474914 655634
rect 474294 619954 474914 655398
rect 474294 619718 474326 619954
rect 474562 619718 474646 619954
rect 474882 619718 474914 619954
rect 474294 619634 474914 619718
rect 474294 619398 474326 619634
rect 474562 619398 474646 619634
rect 474882 619398 474914 619634
rect 380272 583954 380620 583986
rect 380272 583718 380328 583954
rect 380564 583718 380620 583954
rect 380272 583634 380620 583718
rect 380272 583398 380328 583634
rect 380564 583398 380620 583634
rect 380272 583366 380620 583398
rect 470440 583954 470788 583986
rect 470440 583718 470496 583954
rect 470732 583718 470788 583954
rect 470440 583634 470788 583718
rect 470440 583398 470496 583634
rect 470732 583398 470788 583634
rect 470440 583366 470788 583398
rect 474294 583954 474914 619398
rect 474294 583718 474326 583954
rect 474562 583718 474646 583954
rect 474882 583718 474914 583954
rect 474294 583634 474914 583718
rect 474294 583398 474326 583634
rect 474562 583398 474646 583634
rect 474882 583398 474914 583634
rect 380952 579454 381300 579486
rect 380952 579218 381008 579454
rect 381244 579218 381300 579454
rect 380952 579134 381300 579218
rect 380952 578898 381008 579134
rect 381244 578898 381300 579134
rect 380952 578866 381300 578898
rect 469760 579454 470108 579486
rect 469760 579218 469816 579454
rect 470052 579218 470108 579454
rect 469760 579134 470108 579218
rect 469760 578898 469816 579134
rect 470052 578898 470108 579134
rect 469760 578866 470108 578898
rect 375294 556718 375326 556954
rect 375562 556718 375646 556954
rect 375882 556718 375914 556954
rect 375294 556634 375914 556718
rect 375294 556398 375326 556634
rect 375562 556398 375646 556634
rect 375882 556398 375914 556634
rect 375294 520954 375914 556398
rect 380272 547954 380620 547986
rect 380272 547718 380328 547954
rect 380564 547718 380620 547954
rect 380272 547634 380620 547718
rect 380272 547398 380328 547634
rect 380564 547398 380620 547634
rect 380272 547366 380620 547398
rect 470440 547954 470788 547986
rect 470440 547718 470496 547954
rect 470732 547718 470788 547954
rect 470440 547634 470788 547718
rect 470440 547398 470496 547634
rect 470732 547398 470788 547634
rect 470440 547366 470788 547398
rect 474294 547954 474914 583398
rect 474294 547718 474326 547954
rect 474562 547718 474646 547954
rect 474882 547718 474914 547954
rect 474294 547634 474914 547718
rect 474294 547398 474326 547634
rect 474562 547398 474646 547634
rect 474882 547398 474914 547634
rect 380952 543454 381300 543486
rect 380952 543218 381008 543454
rect 381244 543218 381300 543454
rect 380952 543134 381300 543218
rect 380952 542898 381008 543134
rect 381244 542898 381300 543134
rect 380952 542866 381300 542898
rect 469760 543454 470108 543486
rect 469760 543218 469816 543454
rect 470052 543218 470108 543454
rect 469760 543134 470108 543218
rect 469760 542898 469816 543134
rect 470052 542898 470108 543134
rect 469760 542866 470108 542898
rect 375294 520718 375326 520954
rect 375562 520718 375646 520954
rect 375882 520718 375914 520954
rect 375294 520634 375914 520718
rect 375294 520398 375326 520634
rect 375562 520398 375646 520634
rect 375882 520398 375914 520634
rect 375294 484954 375914 520398
rect 380272 511954 380620 511986
rect 380272 511718 380328 511954
rect 380564 511718 380620 511954
rect 380272 511634 380620 511718
rect 380272 511398 380328 511634
rect 380564 511398 380620 511634
rect 380272 511366 380620 511398
rect 470440 511954 470788 511986
rect 470440 511718 470496 511954
rect 470732 511718 470788 511954
rect 470440 511634 470788 511718
rect 470440 511398 470496 511634
rect 470732 511398 470788 511634
rect 470440 511366 470788 511398
rect 474294 511954 474914 547398
rect 474294 511718 474326 511954
rect 474562 511718 474646 511954
rect 474882 511718 474914 511954
rect 474294 511634 474914 511718
rect 474294 511398 474326 511634
rect 474562 511398 474646 511634
rect 474882 511398 474914 511634
rect 380952 507454 381300 507486
rect 380952 507218 381008 507454
rect 381244 507218 381300 507454
rect 380952 507134 381300 507218
rect 380952 506898 381008 507134
rect 381244 506898 381300 507134
rect 380952 506866 381300 506898
rect 469760 507454 470108 507486
rect 469760 507218 469816 507454
rect 470052 507218 470108 507454
rect 469760 507134 470108 507218
rect 469760 506898 469816 507134
rect 470052 506898 470108 507134
rect 469760 506866 470108 506898
rect 392928 499590 392988 500106
rect 394288 499590 394348 500106
rect 395376 499590 395436 500106
rect 397688 499590 397748 500106
rect 392902 499530 392988 499590
rect 394190 499530 394348 499590
rect 395294 499530 395436 499590
rect 397686 499530 397748 499590
rect 398912 499590 398972 500106
rect 400000 499590 400060 500106
rect 401088 499590 401148 500106
rect 402312 499590 402372 500106
rect 403400 499590 403460 500106
rect 404760 499590 404820 500106
rect 405304 499590 405364 500106
rect 398912 499530 399034 499590
rect 375294 484718 375326 484954
rect 375562 484718 375646 484954
rect 375882 484718 375914 484954
rect 375294 484634 375914 484718
rect 375294 484398 375326 484634
rect 375562 484398 375646 484634
rect 375882 484398 375914 484634
rect 375294 448954 375914 484398
rect 375294 448718 375326 448954
rect 375562 448718 375646 448954
rect 375882 448718 375914 448954
rect 375294 448634 375914 448718
rect 375294 448398 375326 448634
rect 375562 448398 375646 448634
rect 375882 448398 375914 448634
rect 375294 412954 375914 448398
rect 375294 412718 375326 412954
rect 375562 412718 375646 412954
rect 375882 412718 375914 412954
rect 375294 412634 375914 412718
rect 375294 412398 375326 412634
rect 375562 412398 375646 412634
rect 375882 412398 375914 412634
rect 375294 376954 375914 412398
rect 375294 376718 375326 376954
rect 375562 376718 375646 376954
rect 375882 376718 375914 376954
rect 375294 376634 375914 376718
rect 375294 376398 375326 376634
rect 375562 376398 375646 376634
rect 375882 376398 375914 376634
rect 375294 340954 375914 376398
rect 375294 340718 375326 340954
rect 375562 340718 375646 340954
rect 375882 340718 375914 340954
rect 375294 340634 375914 340718
rect 375294 340398 375326 340634
rect 375562 340398 375646 340634
rect 375882 340398 375914 340634
rect 375294 304954 375914 340398
rect 375294 304718 375326 304954
rect 375562 304718 375646 304954
rect 375882 304718 375914 304954
rect 375294 304634 375914 304718
rect 375294 304398 375326 304634
rect 375562 304398 375646 304634
rect 375882 304398 375914 304634
rect 375294 268954 375914 304398
rect 375294 268718 375326 268954
rect 375562 268718 375646 268954
rect 375882 268718 375914 268954
rect 375294 268634 375914 268718
rect 375294 268398 375326 268634
rect 375562 268398 375646 268634
rect 375882 268398 375914 268634
rect 375294 232954 375914 268398
rect 375294 232718 375326 232954
rect 375562 232718 375646 232954
rect 375882 232718 375914 232954
rect 375294 232634 375914 232718
rect 375294 232398 375326 232634
rect 375562 232398 375646 232634
rect 375882 232398 375914 232634
rect 375294 196954 375914 232398
rect 375294 196718 375326 196954
rect 375562 196718 375646 196954
rect 375882 196718 375914 196954
rect 375294 196634 375914 196718
rect 375294 196398 375326 196634
rect 375562 196398 375646 196634
rect 375882 196398 375914 196634
rect 375294 160954 375914 196398
rect 375294 160718 375326 160954
rect 375562 160718 375646 160954
rect 375882 160718 375914 160954
rect 375294 160634 375914 160718
rect 375294 160398 375326 160634
rect 375562 160398 375646 160634
rect 375882 160398 375914 160634
rect 375294 124954 375914 160398
rect 375294 124718 375326 124954
rect 375562 124718 375646 124954
rect 375882 124718 375914 124954
rect 375294 124634 375914 124718
rect 375294 124398 375326 124634
rect 375562 124398 375646 124634
rect 375882 124398 375914 124634
rect 375294 88954 375914 124398
rect 375294 88718 375326 88954
rect 375562 88718 375646 88954
rect 375882 88718 375914 88954
rect 375294 88634 375914 88718
rect 375294 88398 375326 88634
rect 375562 88398 375646 88634
rect 375882 88398 375914 88634
rect 375294 52954 375914 88398
rect 375294 52718 375326 52954
rect 375562 52718 375646 52954
rect 375882 52718 375914 52954
rect 375294 52634 375914 52718
rect 375294 52398 375326 52634
rect 375562 52398 375646 52634
rect 375882 52398 375914 52634
rect 375294 16954 375914 52398
rect 375294 16718 375326 16954
rect 375562 16718 375646 16954
rect 375882 16718 375914 16954
rect 375294 16634 375914 16718
rect 375294 16398 375326 16634
rect 375562 16398 375646 16634
rect 375882 16398 375914 16634
rect 375294 -3226 375914 16398
rect 375294 -3462 375326 -3226
rect 375562 -3462 375646 -3226
rect 375882 -3462 375914 -3226
rect 375294 -3546 375914 -3462
rect 375294 -3782 375326 -3546
rect 375562 -3782 375646 -3546
rect 375882 -3782 375914 -3546
rect 375294 -7654 375914 -3782
rect 379794 489454 380414 498000
rect 379794 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 380414 489454
rect 379794 489134 380414 489218
rect 379794 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 380414 489134
rect 379794 453454 380414 488898
rect 379794 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 380414 453454
rect 379794 453134 380414 453218
rect 379794 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 380414 453134
rect 379794 417454 380414 452898
rect 379794 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 380414 417454
rect 379794 417134 380414 417218
rect 379794 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 380414 417134
rect 379794 381454 380414 416898
rect 379794 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 380414 381454
rect 379794 381134 380414 381218
rect 379794 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 380414 381134
rect 379794 345454 380414 380898
rect 379794 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 380414 345454
rect 379794 345134 380414 345218
rect 379794 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 380414 345134
rect 379794 309454 380414 344898
rect 379794 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 380414 309454
rect 379794 309134 380414 309218
rect 379794 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 380414 309134
rect 379794 273454 380414 308898
rect 379794 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 380414 273454
rect 379794 273134 380414 273218
rect 379794 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 380414 273134
rect 379794 237454 380414 272898
rect 379794 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 380414 237454
rect 379794 237134 380414 237218
rect 379794 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 380414 237134
rect 379794 201454 380414 236898
rect 379794 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 380414 201454
rect 379794 201134 380414 201218
rect 379794 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 380414 201134
rect 379794 165454 380414 200898
rect 379794 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 380414 165454
rect 379794 165134 380414 165218
rect 379794 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 380414 165134
rect 379794 129454 380414 164898
rect 379794 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 380414 129454
rect 379794 129134 380414 129218
rect 379794 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 380414 129134
rect 379794 93454 380414 128898
rect 379794 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 380414 93454
rect 379794 93134 380414 93218
rect 379794 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 380414 93134
rect 379794 57454 380414 92898
rect 379794 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 380414 57454
rect 379794 57134 380414 57218
rect 379794 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 380414 57134
rect 379794 21454 380414 56898
rect 379794 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 380414 21454
rect 379794 21134 380414 21218
rect 379794 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 380414 21134
rect 379794 -4186 380414 20898
rect 379794 -4422 379826 -4186
rect 380062 -4422 380146 -4186
rect 380382 -4422 380414 -4186
rect 379794 -4506 380414 -4422
rect 379794 -4742 379826 -4506
rect 380062 -4742 380146 -4506
rect 380382 -4742 380414 -4506
rect 379794 -7654 380414 -4742
rect 384294 493954 384914 498000
rect 384294 493718 384326 493954
rect 384562 493718 384646 493954
rect 384882 493718 384914 493954
rect 384294 493634 384914 493718
rect 384294 493398 384326 493634
rect 384562 493398 384646 493634
rect 384882 493398 384914 493634
rect 384294 457954 384914 493398
rect 384294 457718 384326 457954
rect 384562 457718 384646 457954
rect 384882 457718 384914 457954
rect 384294 457634 384914 457718
rect 384294 457398 384326 457634
rect 384562 457398 384646 457634
rect 384882 457398 384914 457634
rect 384294 421954 384914 457398
rect 384294 421718 384326 421954
rect 384562 421718 384646 421954
rect 384882 421718 384914 421954
rect 384294 421634 384914 421718
rect 384294 421398 384326 421634
rect 384562 421398 384646 421634
rect 384882 421398 384914 421634
rect 384294 385954 384914 421398
rect 384294 385718 384326 385954
rect 384562 385718 384646 385954
rect 384882 385718 384914 385954
rect 384294 385634 384914 385718
rect 384294 385398 384326 385634
rect 384562 385398 384646 385634
rect 384882 385398 384914 385634
rect 384294 349954 384914 385398
rect 384294 349718 384326 349954
rect 384562 349718 384646 349954
rect 384882 349718 384914 349954
rect 384294 349634 384914 349718
rect 384294 349398 384326 349634
rect 384562 349398 384646 349634
rect 384882 349398 384914 349634
rect 384294 313954 384914 349398
rect 384294 313718 384326 313954
rect 384562 313718 384646 313954
rect 384882 313718 384914 313954
rect 384294 313634 384914 313718
rect 384294 313398 384326 313634
rect 384562 313398 384646 313634
rect 384882 313398 384914 313634
rect 384294 277954 384914 313398
rect 384294 277718 384326 277954
rect 384562 277718 384646 277954
rect 384882 277718 384914 277954
rect 384294 277634 384914 277718
rect 384294 277398 384326 277634
rect 384562 277398 384646 277634
rect 384882 277398 384914 277634
rect 384294 241954 384914 277398
rect 384294 241718 384326 241954
rect 384562 241718 384646 241954
rect 384882 241718 384914 241954
rect 384294 241634 384914 241718
rect 384294 241398 384326 241634
rect 384562 241398 384646 241634
rect 384882 241398 384914 241634
rect 384294 205954 384914 241398
rect 384294 205718 384326 205954
rect 384562 205718 384646 205954
rect 384882 205718 384914 205954
rect 384294 205634 384914 205718
rect 384294 205398 384326 205634
rect 384562 205398 384646 205634
rect 384882 205398 384914 205634
rect 384294 169954 384914 205398
rect 384294 169718 384326 169954
rect 384562 169718 384646 169954
rect 384882 169718 384914 169954
rect 384294 169634 384914 169718
rect 384294 169398 384326 169634
rect 384562 169398 384646 169634
rect 384882 169398 384914 169634
rect 384294 133954 384914 169398
rect 384294 133718 384326 133954
rect 384562 133718 384646 133954
rect 384882 133718 384914 133954
rect 384294 133634 384914 133718
rect 384294 133398 384326 133634
rect 384562 133398 384646 133634
rect 384882 133398 384914 133634
rect 384294 97954 384914 133398
rect 384294 97718 384326 97954
rect 384562 97718 384646 97954
rect 384882 97718 384914 97954
rect 384294 97634 384914 97718
rect 384294 97398 384326 97634
rect 384562 97398 384646 97634
rect 384882 97398 384914 97634
rect 384294 61954 384914 97398
rect 384294 61718 384326 61954
rect 384562 61718 384646 61954
rect 384882 61718 384914 61954
rect 384294 61634 384914 61718
rect 384294 61398 384326 61634
rect 384562 61398 384646 61634
rect 384882 61398 384914 61634
rect 384294 25954 384914 61398
rect 384294 25718 384326 25954
rect 384562 25718 384646 25954
rect 384882 25718 384914 25954
rect 384294 25634 384914 25718
rect 384294 25398 384326 25634
rect 384562 25398 384646 25634
rect 384882 25398 384914 25634
rect 384294 -5146 384914 25398
rect 384294 -5382 384326 -5146
rect 384562 -5382 384646 -5146
rect 384882 -5382 384914 -5146
rect 384294 -5466 384914 -5382
rect 384294 -5702 384326 -5466
rect 384562 -5702 384646 -5466
rect 384882 -5702 384914 -5466
rect 384294 -7654 384914 -5702
rect 388794 462454 389414 498000
rect 392902 496909 392962 499530
rect 392899 496908 392965 496909
rect 392899 496844 392900 496908
rect 392964 496844 392965 496908
rect 392899 496843 392965 496844
rect 388794 462218 388826 462454
rect 389062 462218 389146 462454
rect 389382 462218 389414 462454
rect 388794 462134 389414 462218
rect 388794 461898 388826 462134
rect 389062 461898 389146 462134
rect 389382 461898 389414 462134
rect 388794 426454 389414 461898
rect 388794 426218 388826 426454
rect 389062 426218 389146 426454
rect 389382 426218 389414 426454
rect 388794 426134 389414 426218
rect 388794 425898 388826 426134
rect 389062 425898 389146 426134
rect 389382 425898 389414 426134
rect 388794 390454 389414 425898
rect 388794 390218 388826 390454
rect 389062 390218 389146 390454
rect 389382 390218 389414 390454
rect 388794 390134 389414 390218
rect 388794 389898 388826 390134
rect 389062 389898 389146 390134
rect 389382 389898 389414 390134
rect 388794 354454 389414 389898
rect 388794 354218 388826 354454
rect 389062 354218 389146 354454
rect 389382 354218 389414 354454
rect 388794 354134 389414 354218
rect 388794 353898 388826 354134
rect 389062 353898 389146 354134
rect 389382 353898 389414 354134
rect 388794 318454 389414 353898
rect 388794 318218 388826 318454
rect 389062 318218 389146 318454
rect 389382 318218 389414 318454
rect 388794 318134 389414 318218
rect 388794 317898 388826 318134
rect 389062 317898 389146 318134
rect 389382 317898 389414 318134
rect 388794 282454 389414 317898
rect 388794 282218 388826 282454
rect 389062 282218 389146 282454
rect 389382 282218 389414 282454
rect 388794 282134 389414 282218
rect 388794 281898 388826 282134
rect 389062 281898 389146 282134
rect 389382 281898 389414 282134
rect 388794 246454 389414 281898
rect 388794 246218 388826 246454
rect 389062 246218 389146 246454
rect 389382 246218 389414 246454
rect 388794 246134 389414 246218
rect 388794 245898 388826 246134
rect 389062 245898 389146 246134
rect 389382 245898 389414 246134
rect 388794 210454 389414 245898
rect 388794 210218 388826 210454
rect 389062 210218 389146 210454
rect 389382 210218 389414 210454
rect 388794 210134 389414 210218
rect 388794 209898 388826 210134
rect 389062 209898 389146 210134
rect 389382 209898 389414 210134
rect 388794 174454 389414 209898
rect 388794 174218 388826 174454
rect 389062 174218 389146 174454
rect 389382 174218 389414 174454
rect 388794 174134 389414 174218
rect 388794 173898 388826 174134
rect 389062 173898 389146 174134
rect 389382 173898 389414 174134
rect 388794 138454 389414 173898
rect 388794 138218 388826 138454
rect 389062 138218 389146 138454
rect 389382 138218 389414 138454
rect 388794 138134 389414 138218
rect 388794 137898 388826 138134
rect 389062 137898 389146 138134
rect 389382 137898 389414 138134
rect 388794 102454 389414 137898
rect 388794 102218 388826 102454
rect 389062 102218 389146 102454
rect 389382 102218 389414 102454
rect 388794 102134 389414 102218
rect 388794 101898 388826 102134
rect 389062 101898 389146 102134
rect 389382 101898 389414 102134
rect 388794 66454 389414 101898
rect 388794 66218 388826 66454
rect 389062 66218 389146 66454
rect 389382 66218 389414 66454
rect 388794 66134 389414 66218
rect 388794 65898 388826 66134
rect 389062 65898 389146 66134
rect 389382 65898 389414 66134
rect 388794 30454 389414 65898
rect 388794 30218 388826 30454
rect 389062 30218 389146 30454
rect 389382 30218 389414 30454
rect 388794 30134 389414 30218
rect 388794 29898 388826 30134
rect 389062 29898 389146 30134
rect 389382 29898 389414 30134
rect 388794 -6106 389414 29898
rect 388794 -6342 388826 -6106
rect 389062 -6342 389146 -6106
rect 389382 -6342 389414 -6106
rect 388794 -6426 389414 -6342
rect 388794 -6662 388826 -6426
rect 389062 -6662 389146 -6426
rect 389382 -6662 389414 -6426
rect 388794 -7654 389414 -6662
rect 393294 466954 393914 498000
rect 394190 496909 394250 499530
rect 395294 496909 395354 499530
rect 397686 498133 397746 499530
rect 397683 498132 397749 498133
rect 397683 498068 397684 498132
rect 397748 498068 397749 498132
rect 397683 498067 397749 498068
rect 394187 496908 394253 496909
rect 394187 496844 394188 496908
rect 394252 496844 394253 496908
rect 394187 496843 394253 496844
rect 395291 496908 395357 496909
rect 395291 496844 395292 496908
rect 395356 496844 395357 496908
rect 395291 496843 395357 496844
rect 393294 466718 393326 466954
rect 393562 466718 393646 466954
rect 393882 466718 393914 466954
rect 393294 466634 393914 466718
rect 393294 466398 393326 466634
rect 393562 466398 393646 466634
rect 393882 466398 393914 466634
rect 393294 430954 393914 466398
rect 393294 430718 393326 430954
rect 393562 430718 393646 430954
rect 393882 430718 393914 430954
rect 393294 430634 393914 430718
rect 393294 430398 393326 430634
rect 393562 430398 393646 430634
rect 393882 430398 393914 430634
rect 393294 394954 393914 430398
rect 393294 394718 393326 394954
rect 393562 394718 393646 394954
rect 393882 394718 393914 394954
rect 393294 394634 393914 394718
rect 393294 394398 393326 394634
rect 393562 394398 393646 394634
rect 393882 394398 393914 394634
rect 393294 358954 393914 394398
rect 393294 358718 393326 358954
rect 393562 358718 393646 358954
rect 393882 358718 393914 358954
rect 393294 358634 393914 358718
rect 393294 358398 393326 358634
rect 393562 358398 393646 358634
rect 393882 358398 393914 358634
rect 393294 322954 393914 358398
rect 393294 322718 393326 322954
rect 393562 322718 393646 322954
rect 393882 322718 393914 322954
rect 393294 322634 393914 322718
rect 393294 322398 393326 322634
rect 393562 322398 393646 322634
rect 393882 322398 393914 322634
rect 393294 286954 393914 322398
rect 393294 286718 393326 286954
rect 393562 286718 393646 286954
rect 393882 286718 393914 286954
rect 393294 286634 393914 286718
rect 393294 286398 393326 286634
rect 393562 286398 393646 286634
rect 393882 286398 393914 286634
rect 393294 250954 393914 286398
rect 393294 250718 393326 250954
rect 393562 250718 393646 250954
rect 393882 250718 393914 250954
rect 393294 250634 393914 250718
rect 393294 250398 393326 250634
rect 393562 250398 393646 250634
rect 393882 250398 393914 250634
rect 393294 214954 393914 250398
rect 393294 214718 393326 214954
rect 393562 214718 393646 214954
rect 393882 214718 393914 214954
rect 393294 214634 393914 214718
rect 393294 214398 393326 214634
rect 393562 214398 393646 214634
rect 393882 214398 393914 214634
rect 393294 178954 393914 214398
rect 393294 178718 393326 178954
rect 393562 178718 393646 178954
rect 393882 178718 393914 178954
rect 393294 178634 393914 178718
rect 393294 178398 393326 178634
rect 393562 178398 393646 178634
rect 393882 178398 393914 178634
rect 393294 142954 393914 178398
rect 393294 142718 393326 142954
rect 393562 142718 393646 142954
rect 393882 142718 393914 142954
rect 393294 142634 393914 142718
rect 393294 142398 393326 142634
rect 393562 142398 393646 142634
rect 393882 142398 393914 142634
rect 393294 106954 393914 142398
rect 393294 106718 393326 106954
rect 393562 106718 393646 106954
rect 393882 106718 393914 106954
rect 393294 106634 393914 106718
rect 393294 106398 393326 106634
rect 393562 106398 393646 106634
rect 393882 106398 393914 106634
rect 393294 70954 393914 106398
rect 393294 70718 393326 70954
rect 393562 70718 393646 70954
rect 393882 70718 393914 70954
rect 393294 70634 393914 70718
rect 393294 70398 393326 70634
rect 393562 70398 393646 70634
rect 393882 70398 393914 70634
rect 393294 34954 393914 70398
rect 393294 34718 393326 34954
rect 393562 34718 393646 34954
rect 393882 34718 393914 34954
rect 393294 34634 393914 34718
rect 393294 34398 393326 34634
rect 393562 34398 393646 34634
rect 393882 34398 393914 34634
rect 393294 -7066 393914 34398
rect 393294 -7302 393326 -7066
rect 393562 -7302 393646 -7066
rect 393882 -7302 393914 -7066
rect 393294 -7386 393914 -7302
rect 393294 -7622 393326 -7386
rect 393562 -7622 393646 -7386
rect 393882 -7622 393914 -7386
rect 393294 -7654 393914 -7622
rect 397794 471454 398414 498000
rect 398974 497181 399034 499530
rect 399894 499530 400060 499590
rect 400998 499530 401148 499590
rect 402102 499530 402372 499590
rect 403390 499530 403460 499590
rect 404678 499530 404820 499590
rect 405230 499530 405364 499590
rect 405712 499590 405772 500106
rect 410472 499590 410532 500106
rect 405712 499530 405842 499590
rect 399894 497317 399954 499530
rect 399891 497316 399957 497317
rect 399891 497252 399892 497316
rect 399956 497252 399957 497316
rect 399891 497251 399957 497252
rect 398971 497180 399037 497181
rect 398971 497116 398972 497180
rect 399036 497116 399037 497180
rect 398971 497115 399037 497116
rect 400998 496909 401058 499530
rect 402102 496909 402162 499530
rect 400995 496908 401061 496909
rect 400995 496844 400996 496908
rect 401060 496844 401061 496908
rect 400995 496843 401061 496844
rect 402099 496908 402165 496909
rect 402099 496844 402100 496908
rect 402164 496844 402165 496908
rect 402099 496843 402165 496844
rect 397794 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 398414 471454
rect 397794 471134 398414 471218
rect 397794 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 398414 471134
rect 397794 435454 398414 470898
rect 397794 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 398414 435454
rect 397794 435134 398414 435218
rect 397794 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 398414 435134
rect 397794 399454 398414 434898
rect 397794 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 398414 399454
rect 397794 399134 398414 399218
rect 397794 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 398414 399134
rect 397794 363454 398414 398898
rect 397794 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 398414 363454
rect 397794 363134 398414 363218
rect 397794 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 398414 363134
rect 397794 327454 398414 362898
rect 397794 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 398414 327454
rect 397794 327134 398414 327218
rect 397794 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 398414 327134
rect 397794 291454 398414 326898
rect 397794 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 398414 291454
rect 397794 291134 398414 291218
rect 397794 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 398414 291134
rect 397794 255454 398414 290898
rect 397794 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 398414 255454
rect 397794 255134 398414 255218
rect 397794 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 398414 255134
rect 397794 219454 398414 254898
rect 397794 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 398414 219454
rect 397794 219134 398414 219218
rect 397794 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 398414 219134
rect 397794 183454 398414 218898
rect 397794 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 398414 183454
rect 397794 183134 398414 183218
rect 397794 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 398414 183134
rect 397794 147454 398414 182898
rect 397794 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 398414 147454
rect 397794 147134 398414 147218
rect 397794 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 398414 147134
rect 397794 111454 398414 146898
rect 397794 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 398414 111454
rect 397794 111134 398414 111218
rect 397794 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 398414 111134
rect 397794 75454 398414 110898
rect 397794 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 398414 75454
rect 397794 75134 398414 75218
rect 397794 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 398414 75134
rect 397794 39454 398414 74898
rect 397794 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 398414 39454
rect 397794 39134 398414 39218
rect 397794 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 398414 39134
rect 397794 3454 398414 38898
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -7654 398414 -902
rect 402294 475954 402914 498000
rect 403390 497317 403450 499530
rect 403387 497316 403453 497317
rect 403387 497252 403388 497316
rect 403452 497252 403453 497316
rect 403387 497251 403453 497252
rect 404678 496909 404738 499530
rect 405230 497045 405290 499530
rect 405227 497044 405293 497045
rect 405227 496980 405228 497044
rect 405292 496980 405293 497044
rect 405227 496979 405293 496980
rect 405782 496909 405842 499530
rect 410382 499530 410532 499590
rect 415504 499590 415564 500106
rect 420536 499590 420596 500106
rect 425568 499590 425628 500106
rect 430464 499590 430524 500106
rect 435496 499590 435556 500106
rect 415504 499530 415594 499590
rect 404675 496908 404741 496909
rect 404675 496844 404676 496908
rect 404740 496844 404741 496908
rect 404675 496843 404741 496844
rect 405779 496908 405845 496909
rect 405779 496844 405780 496908
rect 405844 496844 405845 496908
rect 405779 496843 405845 496844
rect 402294 475718 402326 475954
rect 402562 475718 402646 475954
rect 402882 475718 402914 475954
rect 402294 475634 402914 475718
rect 402294 475398 402326 475634
rect 402562 475398 402646 475634
rect 402882 475398 402914 475634
rect 402294 439954 402914 475398
rect 402294 439718 402326 439954
rect 402562 439718 402646 439954
rect 402882 439718 402914 439954
rect 402294 439634 402914 439718
rect 402294 439398 402326 439634
rect 402562 439398 402646 439634
rect 402882 439398 402914 439634
rect 402294 403954 402914 439398
rect 402294 403718 402326 403954
rect 402562 403718 402646 403954
rect 402882 403718 402914 403954
rect 402294 403634 402914 403718
rect 402294 403398 402326 403634
rect 402562 403398 402646 403634
rect 402882 403398 402914 403634
rect 402294 367954 402914 403398
rect 402294 367718 402326 367954
rect 402562 367718 402646 367954
rect 402882 367718 402914 367954
rect 402294 367634 402914 367718
rect 402294 367398 402326 367634
rect 402562 367398 402646 367634
rect 402882 367398 402914 367634
rect 402294 331954 402914 367398
rect 402294 331718 402326 331954
rect 402562 331718 402646 331954
rect 402882 331718 402914 331954
rect 402294 331634 402914 331718
rect 402294 331398 402326 331634
rect 402562 331398 402646 331634
rect 402882 331398 402914 331634
rect 402294 295954 402914 331398
rect 402294 295718 402326 295954
rect 402562 295718 402646 295954
rect 402882 295718 402914 295954
rect 402294 295634 402914 295718
rect 402294 295398 402326 295634
rect 402562 295398 402646 295634
rect 402882 295398 402914 295634
rect 402294 259954 402914 295398
rect 402294 259718 402326 259954
rect 402562 259718 402646 259954
rect 402882 259718 402914 259954
rect 402294 259634 402914 259718
rect 402294 259398 402326 259634
rect 402562 259398 402646 259634
rect 402882 259398 402914 259634
rect 402294 223954 402914 259398
rect 402294 223718 402326 223954
rect 402562 223718 402646 223954
rect 402882 223718 402914 223954
rect 402294 223634 402914 223718
rect 402294 223398 402326 223634
rect 402562 223398 402646 223634
rect 402882 223398 402914 223634
rect 402294 187954 402914 223398
rect 402294 187718 402326 187954
rect 402562 187718 402646 187954
rect 402882 187718 402914 187954
rect 402294 187634 402914 187718
rect 402294 187398 402326 187634
rect 402562 187398 402646 187634
rect 402882 187398 402914 187634
rect 402294 151954 402914 187398
rect 402294 151718 402326 151954
rect 402562 151718 402646 151954
rect 402882 151718 402914 151954
rect 402294 151634 402914 151718
rect 402294 151398 402326 151634
rect 402562 151398 402646 151634
rect 402882 151398 402914 151634
rect 402294 115954 402914 151398
rect 402294 115718 402326 115954
rect 402562 115718 402646 115954
rect 402882 115718 402914 115954
rect 402294 115634 402914 115718
rect 402294 115398 402326 115634
rect 402562 115398 402646 115634
rect 402882 115398 402914 115634
rect 402294 79954 402914 115398
rect 402294 79718 402326 79954
rect 402562 79718 402646 79954
rect 402882 79718 402914 79954
rect 402294 79634 402914 79718
rect 402294 79398 402326 79634
rect 402562 79398 402646 79634
rect 402882 79398 402914 79634
rect 402294 43954 402914 79398
rect 402294 43718 402326 43954
rect 402562 43718 402646 43954
rect 402882 43718 402914 43954
rect 402294 43634 402914 43718
rect 402294 43398 402326 43634
rect 402562 43398 402646 43634
rect 402882 43398 402914 43634
rect 402294 7954 402914 43398
rect 402294 7718 402326 7954
rect 402562 7718 402646 7954
rect 402882 7718 402914 7954
rect 402294 7634 402914 7718
rect 402294 7398 402326 7634
rect 402562 7398 402646 7634
rect 402882 7398 402914 7634
rect 402294 -1306 402914 7398
rect 402294 -1542 402326 -1306
rect 402562 -1542 402646 -1306
rect 402882 -1542 402914 -1306
rect 402294 -1626 402914 -1542
rect 402294 -1862 402326 -1626
rect 402562 -1862 402646 -1626
rect 402882 -1862 402914 -1626
rect 402294 -7654 402914 -1862
rect 406794 480454 407414 498000
rect 410382 497725 410442 499530
rect 410379 497724 410445 497725
rect 410379 497660 410380 497724
rect 410444 497660 410445 497724
rect 410379 497659 410445 497660
rect 406794 480218 406826 480454
rect 407062 480218 407146 480454
rect 407382 480218 407414 480454
rect 406794 480134 407414 480218
rect 406794 479898 406826 480134
rect 407062 479898 407146 480134
rect 407382 479898 407414 480134
rect 406794 444454 407414 479898
rect 406794 444218 406826 444454
rect 407062 444218 407146 444454
rect 407382 444218 407414 444454
rect 406794 444134 407414 444218
rect 406794 443898 406826 444134
rect 407062 443898 407146 444134
rect 407382 443898 407414 444134
rect 406794 408454 407414 443898
rect 406794 408218 406826 408454
rect 407062 408218 407146 408454
rect 407382 408218 407414 408454
rect 406794 408134 407414 408218
rect 406794 407898 406826 408134
rect 407062 407898 407146 408134
rect 407382 407898 407414 408134
rect 406794 372454 407414 407898
rect 406794 372218 406826 372454
rect 407062 372218 407146 372454
rect 407382 372218 407414 372454
rect 406794 372134 407414 372218
rect 406794 371898 406826 372134
rect 407062 371898 407146 372134
rect 407382 371898 407414 372134
rect 406794 336454 407414 371898
rect 406794 336218 406826 336454
rect 407062 336218 407146 336454
rect 407382 336218 407414 336454
rect 406794 336134 407414 336218
rect 406794 335898 406826 336134
rect 407062 335898 407146 336134
rect 407382 335898 407414 336134
rect 406794 300454 407414 335898
rect 406794 300218 406826 300454
rect 407062 300218 407146 300454
rect 407382 300218 407414 300454
rect 406794 300134 407414 300218
rect 406794 299898 406826 300134
rect 407062 299898 407146 300134
rect 407382 299898 407414 300134
rect 406794 264454 407414 299898
rect 406794 264218 406826 264454
rect 407062 264218 407146 264454
rect 407382 264218 407414 264454
rect 406794 264134 407414 264218
rect 406794 263898 406826 264134
rect 407062 263898 407146 264134
rect 407382 263898 407414 264134
rect 406794 228454 407414 263898
rect 406794 228218 406826 228454
rect 407062 228218 407146 228454
rect 407382 228218 407414 228454
rect 406794 228134 407414 228218
rect 406794 227898 406826 228134
rect 407062 227898 407146 228134
rect 407382 227898 407414 228134
rect 406794 192454 407414 227898
rect 406794 192218 406826 192454
rect 407062 192218 407146 192454
rect 407382 192218 407414 192454
rect 406794 192134 407414 192218
rect 406794 191898 406826 192134
rect 407062 191898 407146 192134
rect 407382 191898 407414 192134
rect 406794 156454 407414 191898
rect 406794 156218 406826 156454
rect 407062 156218 407146 156454
rect 407382 156218 407414 156454
rect 406794 156134 407414 156218
rect 406794 155898 406826 156134
rect 407062 155898 407146 156134
rect 407382 155898 407414 156134
rect 406794 120454 407414 155898
rect 406794 120218 406826 120454
rect 407062 120218 407146 120454
rect 407382 120218 407414 120454
rect 406794 120134 407414 120218
rect 406794 119898 406826 120134
rect 407062 119898 407146 120134
rect 407382 119898 407414 120134
rect 406794 84454 407414 119898
rect 406794 84218 406826 84454
rect 407062 84218 407146 84454
rect 407382 84218 407414 84454
rect 406794 84134 407414 84218
rect 406794 83898 406826 84134
rect 407062 83898 407146 84134
rect 407382 83898 407414 84134
rect 406794 48454 407414 83898
rect 406794 48218 406826 48454
rect 407062 48218 407146 48454
rect 407382 48218 407414 48454
rect 406794 48134 407414 48218
rect 406794 47898 406826 48134
rect 407062 47898 407146 48134
rect 407382 47898 407414 48134
rect 406794 12454 407414 47898
rect 406794 12218 406826 12454
rect 407062 12218 407146 12454
rect 407382 12218 407414 12454
rect 406794 12134 407414 12218
rect 406794 11898 406826 12134
rect 407062 11898 407146 12134
rect 407382 11898 407414 12134
rect 406794 -2266 407414 11898
rect 406794 -2502 406826 -2266
rect 407062 -2502 407146 -2266
rect 407382 -2502 407414 -2266
rect 406794 -2586 407414 -2502
rect 406794 -2822 406826 -2586
rect 407062 -2822 407146 -2586
rect 407382 -2822 407414 -2586
rect 406794 -7654 407414 -2822
rect 411294 484954 411914 498000
rect 415534 496909 415594 499530
rect 420134 499530 420596 499590
rect 425470 499530 425628 499590
rect 430438 499530 430524 499590
rect 435406 499530 435556 499590
rect 440528 499590 440588 500106
rect 440528 499530 440618 499590
rect 415531 496908 415597 496909
rect 415531 496844 415532 496908
rect 415596 496844 415597 496908
rect 415531 496843 415597 496844
rect 411294 484718 411326 484954
rect 411562 484718 411646 484954
rect 411882 484718 411914 484954
rect 411294 484634 411914 484718
rect 411294 484398 411326 484634
rect 411562 484398 411646 484634
rect 411882 484398 411914 484634
rect 411294 448954 411914 484398
rect 411294 448718 411326 448954
rect 411562 448718 411646 448954
rect 411882 448718 411914 448954
rect 411294 448634 411914 448718
rect 411294 448398 411326 448634
rect 411562 448398 411646 448634
rect 411882 448398 411914 448634
rect 411294 412954 411914 448398
rect 411294 412718 411326 412954
rect 411562 412718 411646 412954
rect 411882 412718 411914 412954
rect 411294 412634 411914 412718
rect 411294 412398 411326 412634
rect 411562 412398 411646 412634
rect 411882 412398 411914 412634
rect 411294 376954 411914 412398
rect 411294 376718 411326 376954
rect 411562 376718 411646 376954
rect 411882 376718 411914 376954
rect 411294 376634 411914 376718
rect 411294 376398 411326 376634
rect 411562 376398 411646 376634
rect 411882 376398 411914 376634
rect 411294 340954 411914 376398
rect 411294 340718 411326 340954
rect 411562 340718 411646 340954
rect 411882 340718 411914 340954
rect 411294 340634 411914 340718
rect 411294 340398 411326 340634
rect 411562 340398 411646 340634
rect 411882 340398 411914 340634
rect 411294 304954 411914 340398
rect 411294 304718 411326 304954
rect 411562 304718 411646 304954
rect 411882 304718 411914 304954
rect 411294 304634 411914 304718
rect 411294 304398 411326 304634
rect 411562 304398 411646 304634
rect 411882 304398 411914 304634
rect 411294 268954 411914 304398
rect 411294 268718 411326 268954
rect 411562 268718 411646 268954
rect 411882 268718 411914 268954
rect 411294 268634 411914 268718
rect 411294 268398 411326 268634
rect 411562 268398 411646 268634
rect 411882 268398 411914 268634
rect 411294 232954 411914 268398
rect 411294 232718 411326 232954
rect 411562 232718 411646 232954
rect 411882 232718 411914 232954
rect 411294 232634 411914 232718
rect 411294 232398 411326 232634
rect 411562 232398 411646 232634
rect 411882 232398 411914 232634
rect 411294 196954 411914 232398
rect 411294 196718 411326 196954
rect 411562 196718 411646 196954
rect 411882 196718 411914 196954
rect 411294 196634 411914 196718
rect 411294 196398 411326 196634
rect 411562 196398 411646 196634
rect 411882 196398 411914 196634
rect 411294 160954 411914 196398
rect 411294 160718 411326 160954
rect 411562 160718 411646 160954
rect 411882 160718 411914 160954
rect 411294 160634 411914 160718
rect 411294 160398 411326 160634
rect 411562 160398 411646 160634
rect 411882 160398 411914 160634
rect 411294 124954 411914 160398
rect 411294 124718 411326 124954
rect 411562 124718 411646 124954
rect 411882 124718 411914 124954
rect 411294 124634 411914 124718
rect 411294 124398 411326 124634
rect 411562 124398 411646 124634
rect 411882 124398 411914 124634
rect 411294 88954 411914 124398
rect 411294 88718 411326 88954
rect 411562 88718 411646 88954
rect 411882 88718 411914 88954
rect 411294 88634 411914 88718
rect 411294 88398 411326 88634
rect 411562 88398 411646 88634
rect 411882 88398 411914 88634
rect 411294 52954 411914 88398
rect 411294 52718 411326 52954
rect 411562 52718 411646 52954
rect 411882 52718 411914 52954
rect 411294 52634 411914 52718
rect 411294 52398 411326 52634
rect 411562 52398 411646 52634
rect 411882 52398 411914 52634
rect 411294 16954 411914 52398
rect 411294 16718 411326 16954
rect 411562 16718 411646 16954
rect 411882 16718 411914 16954
rect 411294 16634 411914 16718
rect 411294 16398 411326 16634
rect 411562 16398 411646 16634
rect 411882 16398 411914 16634
rect 411294 -3226 411914 16398
rect 411294 -3462 411326 -3226
rect 411562 -3462 411646 -3226
rect 411882 -3462 411914 -3226
rect 411294 -3546 411914 -3462
rect 411294 -3782 411326 -3546
rect 411562 -3782 411646 -3546
rect 411882 -3782 411914 -3546
rect 411294 -7654 411914 -3782
rect 415794 489454 416414 498000
rect 420134 496909 420194 499530
rect 425470 498133 425530 499530
rect 425467 498132 425533 498133
rect 425467 498068 425468 498132
rect 425532 498068 425533 498132
rect 425467 498067 425533 498068
rect 420131 496908 420197 496909
rect 420131 496844 420132 496908
rect 420196 496844 420197 496908
rect 420131 496843 420197 496844
rect 415794 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 416414 489454
rect 415794 489134 416414 489218
rect 415794 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 416414 489134
rect 415794 453454 416414 488898
rect 415794 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 416414 453454
rect 415794 453134 416414 453218
rect 415794 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 416414 453134
rect 415794 417454 416414 452898
rect 415794 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 416414 417454
rect 415794 417134 416414 417218
rect 415794 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 416414 417134
rect 415794 381454 416414 416898
rect 415794 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 416414 381454
rect 415794 381134 416414 381218
rect 415794 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 416414 381134
rect 415794 345454 416414 380898
rect 415794 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 416414 345454
rect 415794 345134 416414 345218
rect 415794 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 416414 345134
rect 415794 309454 416414 344898
rect 415794 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 416414 309454
rect 415794 309134 416414 309218
rect 415794 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 416414 309134
rect 415794 273454 416414 308898
rect 415794 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 416414 273454
rect 415794 273134 416414 273218
rect 415794 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 416414 273134
rect 415794 237454 416414 272898
rect 415794 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 416414 237454
rect 415794 237134 416414 237218
rect 415794 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 416414 237134
rect 415794 201454 416414 236898
rect 415794 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 416414 201454
rect 415794 201134 416414 201218
rect 415794 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 416414 201134
rect 415794 165454 416414 200898
rect 415794 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 416414 165454
rect 415794 165134 416414 165218
rect 415794 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 416414 165134
rect 415794 129454 416414 164898
rect 415794 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 416414 129454
rect 415794 129134 416414 129218
rect 415794 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 416414 129134
rect 415794 93454 416414 128898
rect 415794 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 416414 93454
rect 415794 93134 416414 93218
rect 415794 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 416414 93134
rect 415794 57454 416414 92898
rect 415794 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 416414 57454
rect 415794 57134 416414 57218
rect 415794 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 416414 57134
rect 415794 21454 416414 56898
rect 415794 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 416414 21454
rect 415794 21134 416414 21218
rect 415794 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 416414 21134
rect 415794 -4186 416414 20898
rect 415794 -4422 415826 -4186
rect 416062 -4422 416146 -4186
rect 416382 -4422 416414 -4186
rect 415794 -4506 416414 -4422
rect 415794 -4742 415826 -4506
rect 416062 -4742 416146 -4506
rect 416382 -4742 416414 -4506
rect 415794 -7654 416414 -4742
rect 420294 493954 420914 498000
rect 420294 493718 420326 493954
rect 420562 493718 420646 493954
rect 420882 493718 420914 493954
rect 420294 493634 420914 493718
rect 420294 493398 420326 493634
rect 420562 493398 420646 493634
rect 420882 493398 420914 493634
rect 420294 457954 420914 493398
rect 420294 457718 420326 457954
rect 420562 457718 420646 457954
rect 420882 457718 420914 457954
rect 420294 457634 420914 457718
rect 420294 457398 420326 457634
rect 420562 457398 420646 457634
rect 420882 457398 420914 457634
rect 420294 421954 420914 457398
rect 420294 421718 420326 421954
rect 420562 421718 420646 421954
rect 420882 421718 420914 421954
rect 420294 421634 420914 421718
rect 420294 421398 420326 421634
rect 420562 421398 420646 421634
rect 420882 421398 420914 421634
rect 420294 385954 420914 421398
rect 420294 385718 420326 385954
rect 420562 385718 420646 385954
rect 420882 385718 420914 385954
rect 420294 385634 420914 385718
rect 420294 385398 420326 385634
rect 420562 385398 420646 385634
rect 420882 385398 420914 385634
rect 420294 349954 420914 385398
rect 420294 349718 420326 349954
rect 420562 349718 420646 349954
rect 420882 349718 420914 349954
rect 420294 349634 420914 349718
rect 420294 349398 420326 349634
rect 420562 349398 420646 349634
rect 420882 349398 420914 349634
rect 420294 313954 420914 349398
rect 420294 313718 420326 313954
rect 420562 313718 420646 313954
rect 420882 313718 420914 313954
rect 420294 313634 420914 313718
rect 420294 313398 420326 313634
rect 420562 313398 420646 313634
rect 420882 313398 420914 313634
rect 420294 277954 420914 313398
rect 420294 277718 420326 277954
rect 420562 277718 420646 277954
rect 420882 277718 420914 277954
rect 420294 277634 420914 277718
rect 420294 277398 420326 277634
rect 420562 277398 420646 277634
rect 420882 277398 420914 277634
rect 420294 241954 420914 277398
rect 420294 241718 420326 241954
rect 420562 241718 420646 241954
rect 420882 241718 420914 241954
rect 420294 241634 420914 241718
rect 420294 241398 420326 241634
rect 420562 241398 420646 241634
rect 420882 241398 420914 241634
rect 420294 205954 420914 241398
rect 420294 205718 420326 205954
rect 420562 205718 420646 205954
rect 420882 205718 420914 205954
rect 420294 205634 420914 205718
rect 420294 205398 420326 205634
rect 420562 205398 420646 205634
rect 420882 205398 420914 205634
rect 420294 169954 420914 205398
rect 420294 169718 420326 169954
rect 420562 169718 420646 169954
rect 420882 169718 420914 169954
rect 420294 169634 420914 169718
rect 420294 169398 420326 169634
rect 420562 169398 420646 169634
rect 420882 169398 420914 169634
rect 420294 133954 420914 169398
rect 420294 133718 420326 133954
rect 420562 133718 420646 133954
rect 420882 133718 420914 133954
rect 420294 133634 420914 133718
rect 420294 133398 420326 133634
rect 420562 133398 420646 133634
rect 420882 133398 420914 133634
rect 420294 97954 420914 133398
rect 420294 97718 420326 97954
rect 420562 97718 420646 97954
rect 420882 97718 420914 97954
rect 420294 97634 420914 97718
rect 420294 97398 420326 97634
rect 420562 97398 420646 97634
rect 420882 97398 420914 97634
rect 420294 61954 420914 97398
rect 420294 61718 420326 61954
rect 420562 61718 420646 61954
rect 420882 61718 420914 61954
rect 420294 61634 420914 61718
rect 420294 61398 420326 61634
rect 420562 61398 420646 61634
rect 420882 61398 420914 61634
rect 420294 25954 420914 61398
rect 420294 25718 420326 25954
rect 420562 25718 420646 25954
rect 420882 25718 420914 25954
rect 420294 25634 420914 25718
rect 420294 25398 420326 25634
rect 420562 25398 420646 25634
rect 420882 25398 420914 25634
rect 420294 -5146 420914 25398
rect 420294 -5382 420326 -5146
rect 420562 -5382 420646 -5146
rect 420882 -5382 420914 -5146
rect 420294 -5466 420914 -5382
rect 420294 -5702 420326 -5466
rect 420562 -5702 420646 -5466
rect 420882 -5702 420914 -5466
rect 420294 -7654 420914 -5702
rect 424794 462454 425414 498000
rect 424794 462218 424826 462454
rect 425062 462218 425146 462454
rect 425382 462218 425414 462454
rect 424794 462134 425414 462218
rect 424794 461898 424826 462134
rect 425062 461898 425146 462134
rect 425382 461898 425414 462134
rect 424794 426454 425414 461898
rect 424794 426218 424826 426454
rect 425062 426218 425146 426454
rect 425382 426218 425414 426454
rect 424794 426134 425414 426218
rect 424794 425898 424826 426134
rect 425062 425898 425146 426134
rect 425382 425898 425414 426134
rect 424794 390454 425414 425898
rect 424794 390218 424826 390454
rect 425062 390218 425146 390454
rect 425382 390218 425414 390454
rect 424794 390134 425414 390218
rect 424794 389898 424826 390134
rect 425062 389898 425146 390134
rect 425382 389898 425414 390134
rect 424794 354454 425414 389898
rect 424794 354218 424826 354454
rect 425062 354218 425146 354454
rect 425382 354218 425414 354454
rect 424794 354134 425414 354218
rect 424794 353898 424826 354134
rect 425062 353898 425146 354134
rect 425382 353898 425414 354134
rect 424794 318454 425414 353898
rect 424794 318218 424826 318454
rect 425062 318218 425146 318454
rect 425382 318218 425414 318454
rect 424794 318134 425414 318218
rect 424794 317898 424826 318134
rect 425062 317898 425146 318134
rect 425382 317898 425414 318134
rect 424794 282454 425414 317898
rect 424794 282218 424826 282454
rect 425062 282218 425146 282454
rect 425382 282218 425414 282454
rect 424794 282134 425414 282218
rect 424794 281898 424826 282134
rect 425062 281898 425146 282134
rect 425382 281898 425414 282134
rect 424794 246454 425414 281898
rect 424794 246218 424826 246454
rect 425062 246218 425146 246454
rect 425382 246218 425414 246454
rect 424794 246134 425414 246218
rect 424794 245898 424826 246134
rect 425062 245898 425146 246134
rect 425382 245898 425414 246134
rect 424794 210454 425414 245898
rect 424794 210218 424826 210454
rect 425062 210218 425146 210454
rect 425382 210218 425414 210454
rect 424794 210134 425414 210218
rect 424794 209898 424826 210134
rect 425062 209898 425146 210134
rect 425382 209898 425414 210134
rect 424794 174454 425414 209898
rect 424794 174218 424826 174454
rect 425062 174218 425146 174454
rect 425382 174218 425414 174454
rect 424794 174134 425414 174218
rect 424794 173898 424826 174134
rect 425062 173898 425146 174134
rect 425382 173898 425414 174134
rect 424794 138454 425414 173898
rect 424794 138218 424826 138454
rect 425062 138218 425146 138454
rect 425382 138218 425414 138454
rect 424794 138134 425414 138218
rect 424794 137898 424826 138134
rect 425062 137898 425146 138134
rect 425382 137898 425414 138134
rect 424794 102454 425414 137898
rect 424794 102218 424826 102454
rect 425062 102218 425146 102454
rect 425382 102218 425414 102454
rect 424794 102134 425414 102218
rect 424794 101898 424826 102134
rect 425062 101898 425146 102134
rect 425382 101898 425414 102134
rect 424794 66454 425414 101898
rect 424794 66218 424826 66454
rect 425062 66218 425146 66454
rect 425382 66218 425414 66454
rect 424794 66134 425414 66218
rect 424794 65898 424826 66134
rect 425062 65898 425146 66134
rect 425382 65898 425414 66134
rect 424794 30454 425414 65898
rect 424794 30218 424826 30454
rect 425062 30218 425146 30454
rect 425382 30218 425414 30454
rect 424794 30134 425414 30218
rect 424794 29898 424826 30134
rect 425062 29898 425146 30134
rect 425382 29898 425414 30134
rect 424794 -6106 425414 29898
rect 424794 -6342 424826 -6106
rect 425062 -6342 425146 -6106
rect 425382 -6342 425414 -6106
rect 424794 -6426 425414 -6342
rect 424794 -6662 424826 -6426
rect 425062 -6662 425146 -6426
rect 425382 -6662 425414 -6426
rect 424794 -7654 425414 -6662
rect 429294 466954 429914 498000
rect 430438 496909 430498 499530
rect 430435 496908 430501 496909
rect 430435 496844 430436 496908
rect 430500 496844 430501 496908
rect 430435 496843 430501 496844
rect 429294 466718 429326 466954
rect 429562 466718 429646 466954
rect 429882 466718 429914 466954
rect 429294 466634 429914 466718
rect 429294 466398 429326 466634
rect 429562 466398 429646 466634
rect 429882 466398 429914 466634
rect 429294 430954 429914 466398
rect 429294 430718 429326 430954
rect 429562 430718 429646 430954
rect 429882 430718 429914 430954
rect 429294 430634 429914 430718
rect 429294 430398 429326 430634
rect 429562 430398 429646 430634
rect 429882 430398 429914 430634
rect 429294 394954 429914 430398
rect 429294 394718 429326 394954
rect 429562 394718 429646 394954
rect 429882 394718 429914 394954
rect 429294 394634 429914 394718
rect 429294 394398 429326 394634
rect 429562 394398 429646 394634
rect 429882 394398 429914 394634
rect 429294 358954 429914 394398
rect 429294 358718 429326 358954
rect 429562 358718 429646 358954
rect 429882 358718 429914 358954
rect 429294 358634 429914 358718
rect 429294 358398 429326 358634
rect 429562 358398 429646 358634
rect 429882 358398 429914 358634
rect 429294 322954 429914 358398
rect 429294 322718 429326 322954
rect 429562 322718 429646 322954
rect 429882 322718 429914 322954
rect 429294 322634 429914 322718
rect 429294 322398 429326 322634
rect 429562 322398 429646 322634
rect 429882 322398 429914 322634
rect 429294 286954 429914 322398
rect 429294 286718 429326 286954
rect 429562 286718 429646 286954
rect 429882 286718 429914 286954
rect 429294 286634 429914 286718
rect 429294 286398 429326 286634
rect 429562 286398 429646 286634
rect 429882 286398 429914 286634
rect 429294 250954 429914 286398
rect 429294 250718 429326 250954
rect 429562 250718 429646 250954
rect 429882 250718 429914 250954
rect 429294 250634 429914 250718
rect 429294 250398 429326 250634
rect 429562 250398 429646 250634
rect 429882 250398 429914 250634
rect 429294 214954 429914 250398
rect 429294 214718 429326 214954
rect 429562 214718 429646 214954
rect 429882 214718 429914 214954
rect 429294 214634 429914 214718
rect 429294 214398 429326 214634
rect 429562 214398 429646 214634
rect 429882 214398 429914 214634
rect 429294 178954 429914 214398
rect 429294 178718 429326 178954
rect 429562 178718 429646 178954
rect 429882 178718 429914 178954
rect 429294 178634 429914 178718
rect 429294 178398 429326 178634
rect 429562 178398 429646 178634
rect 429882 178398 429914 178634
rect 429294 142954 429914 178398
rect 429294 142718 429326 142954
rect 429562 142718 429646 142954
rect 429882 142718 429914 142954
rect 429294 142634 429914 142718
rect 429294 142398 429326 142634
rect 429562 142398 429646 142634
rect 429882 142398 429914 142634
rect 429294 106954 429914 142398
rect 429294 106718 429326 106954
rect 429562 106718 429646 106954
rect 429882 106718 429914 106954
rect 429294 106634 429914 106718
rect 429294 106398 429326 106634
rect 429562 106398 429646 106634
rect 429882 106398 429914 106634
rect 429294 70954 429914 106398
rect 429294 70718 429326 70954
rect 429562 70718 429646 70954
rect 429882 70718 429914 70954
rect 429294 70634 429914 70718
rect 429294 70398 429326 70634
rect 429562 70398 429646 70634
rect 429882 70398 429914 70634
rect 429294 34954 429914 70398
rect 429294 34718 429326 34954
rect 429562 34718 429646 34954
rect 429882 34718 429914 34954
rect 429294 34634 429914 34718
rect 429294 34398 429326 34634
rect 429562 34398 429646 34634
rect 429882 34398 429914 34634
rect 429294 -7066 429914 34398
rect 429294 -7302 429326 -7066
rect 429562 -7302 429646 -7066
rect 429882 -7302 429914 -7066
rect 429294 -7386 429914 -7302
rect 429294 -7622 429326 -7386
rect 429562 -7622 429646 -7386
rect 429882 -7622 429914 -7386
rect 429294 -7654 429914 -7622
rect 433794 471454 434414 498000
rect 435406 496909 435466 499530
rect 435403 496908 435469 496909
rect 435403 496844 435404 496908
rect 435468 496844 435469 496908
rect 435403 496843 435469 496844
rect 433794 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 434414 471454
rect 433794 471134 434414 471218
rect 433794 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 434414 471134
rect 433794 435454 434414 470898
rect 433794 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 434414 435454
rect 433794 435134 434414 435218
rect 433794 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 434414 435134
rect 433794 399454 434414 434898
rect 433794 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 434414 399454
rect 433794 399134 434414 399218
rect 433794 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 434414 399134
rect 433794 363454 434414 398898
rect 433794 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 434414 363454
rect 433794 363134 434414 363218
rect 433794 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 434414 363134
rect 433794 327454 434414 362898
rect 433794 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 434414 327454
rect 433794 327134 434414 327218
rect 433794 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 434414 327134
rect 433794 291454 434414 326898
rect 433794 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 434414 291454
rect 433794 291134 434414 291218
rect 433794 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 434414 291134
rect 433794 255454 434414 290898
rect 433794 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 434414 255454
rect 433794 255134 434414 255218
rect 433794 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 434414 255134
rect 433794 219454 434414 254898
rect 433794 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 434414 219454
rect 433794 219134 434414 219218
rect 433794 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 434414 219134
rect 433794 183454 434414 218898
rect 433794 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 434414 183454
rect 433794 183134 434414 183218
rect 433794 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 434414 183134
rect 433794 147454 434414 182898
rect 433794 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 434414 147454
rect 433794 147134 434414 147218
rect 433794 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 434414 147134
rect 433794 111454 434414 146898
rect 433794 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 434414 111454
rect 433794 111134 434414 111218
rect 433794 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 434414 111134
rect 433794 75454 434414 110898
rect 433794 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 434414 75454
rect 433794 75134 434414 75218
rect 433794 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 434414 75134
rect 433794 39454 434414 74898
rect 433794 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 434414 39454
rect 433794 39134 434414 39218
rect 433794 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 434414 39134
rect 433794 3454 434414 38898
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -7654 434414 -902
rect 438294 475954 438914 498000
rect 440558 496909 440618 499530
rect 440555 496908 440621 496909
rect 440555 496844 440556 496908
rect 440620 496844 440621 496908
rect 440555 496843 440621 496844
rect 438294 475718 438326 475954
rect 438562 475718 438646 475954
rect 438882 475718 438914 475954
rect 438294 475634 438914 475718
rect 438294 475398 438326 475634
rect 438562 475398 438646 475634
rect 438882 475398 438914 475634
rect 438294 439954 438914 475398
rect 438294 439718 438326 439954
rect 438562 439718 438646 439954
rect 438882 439718 438914 439954
rect 438294 439634 438914 439718
rect 438294 439398 438326 439634
rect 438562 439398 438646 439634
rect 438882 439398 438914 439634
rect 438294 403954 438914 439398
rect 438294 403718 438326 403954
rect 438562 403718 438646 403954
rect 438882 403718 438914 403954
rect 438294 403634 438914 403718
rect 438294 403398 438326 403634
rect 438562 403398 438646 403634
rect 438882 403398 438914 403634
rect 438294 367954 438914 403398
rect 438294 367718 438326 367954
rect 438562 367718 438646 367954
rect 438882 367718 438914 367954
rect 438294 367634 438914 367718
rect 438294 367398 438326 367634
rect 438562 367398 438646 367634
rect 438882 367398 438914 367634
rect 438294 331954 438914 367398
rect 438294 331718 438326 331954
rect 438562 331718 438646 331954
rect 438882 331718 438914 331954
rect 438294 331634 438914 331718
rect 438294 331398 438326 331634
rect 438562 331398 438646 331634
rect 438882 331398 438914 331634
rect 438294 295954 438914 331398
rect 438294 295718 438326 295954
rect 438562 295718 438646 295954
rect 438882 295718 438914 295954
rect 438294 295634 438914 295718
rect 438294 295398 438326 295634
rect 438562 295398 438646 295634
rect 438882 295398 438914 295634
rect 438294 259954 438914 295398
rect 438294 259718 438326 259954
rect 438562 259718 438646 259954
rect 438882 259718 438914 259954
rect 438294 259634 438914 259718
rect 438294 259398 438326 259634
rect 438562 259398 438646 259634
rect 438882 259398 438914 259634
rect 438294 223954 438914 259398
rect 438294 223718 438326 223954
rect 438562 223718 438646 223954
rect 438882 223718 438914 223954
rect 438294 223634 438914 223718
rect 438294 223398 438326 223634
rect 438562 223398 438646 223634
rect 438882 223398 438914 223634
rect 438294 187954 438914 223398
rect 438294 187718 438326 187954
rect 438562 187718 438646 187954
rect 438882 187718 438914 187954
rect 438294 187634 438914 187718
rect 438294 187398 438326 187634
rect 438562 187398 438646 187634
rect 438882 187398 438914 187634
rect 438294 151954 438914 187398
rect 438294 151718 438326 151954
rect 438562 151718 438646 151954
rect 438882 151718 438914 151954
rect 438294 151634 438914 151718
rect 438294 151398 438326 151634
rect 438562 151398 438646 151634
rect 438882 151398 438914 151634
rect 438294 115954 438914 151398
rect 438294 115718 438326 115954
rect 438562 115718 438646 115954
rect 438882 115718 438914 115954
rect 438294 115634 438914 115718
rect 438294 115398 438326 115634
rect 438562 115398 438646 115634
rect 438882 115398 438914 115634
rect 438294 79954 438914 115398
rect 438294 79718 438326 79954
rect 438562 79718 438646 79954
rect 438882 79718 438914 79954
rect 438294 79634 438914 79718
rect 438294 79398 438326 79634
rect 438562 79398 438646 79634
rect 438882 79398 438914 79634
rect 438294 43954 438914 79398
rect 438294 43718 438326 43954
rect 438562 43718 438646 43954
rect 438882 43718 438914 43954
rect 438294 43634 438914 43718
rect 438294 43398 438326 43634
rect 438562 43398 438646 43634
rect 438882 43398 438914 43634
rect 438294 7954 438914 43398
rect 438294 7718 438326 7954
rect 438562 7718 438646 7954
rect 438882 7718 438914 7954
rect 438294 7634 438914 7718
rect 438294 7398 438326 7634
rect 438562 7398 438646 7634
rect 438882 7398 438914 7634
rect 438294 -1306 438914 7398
rect 438294 -1542 438326 -1306
rect 438562 -1542 438646 -1306
rect 438882 -1542 438914 -1306
rect 438294 -1626 438914 -1542
rect 438294 -1862 438326 -1626
rect 438562 -1862 438646 -1626
rect 438882 -1862 438914 -1626
rect 438294 -7654 438914 -1862
rect 442794 480454 443414 498000
rect 442794 480218 442826 480454
rect 443062 480218 443146 480454
rect 443382 480218 443414 480454
rect 442794 480134 443414 480218
rect 442794 479898 442826 480134
rect 443062 479898 443146 480134
rect 443382 479898 443414 480134
rect 442794 444454 443414 479898
rect 442794 444218 442826 444454
rect 443062 444218 443146 444454
rect 443382 444218 443414 444454
rect 442794 444134 443414 444218
rect 442794 443898 442826 444134
rect 443062 443898 443146 444134
rect 443382 443898 443414 444134
rect 442794 408454 443414 443898
rect 442794 408218 442826 408454
rect 443062 408218 443146 408454
rect 443382 408218 443414 408454
rect 442794 408134 443414 408218
rect 442794 407898 442826 408134
rect 443062 407898 443146 408134
rect 443382 407898 443414 408134
rect 442794 372454 443414 407898
rect 442794 372218 442826 372454
rect 443062 372218 443146 372454
rect 443382 372218 443414 372454
rect 442794 372134 443414 372218
rect 442794 371898 442826 372134
rect 443062 371898 443146 372134
rect 443382 371898 443414 372134
rect 442794 336454 443414 371898
rect 442794 336218 442826 336454
rect 443062 336218 443146 336454
rect 443382 336218 443414 336454
rect 442794 336134 443414 336218
rect 442794 335898 442826 336134
rect 443062 335898 443146 336134
rect 443382 335898 443414 336134
rect 442794 300454 443414 335898
rect 442794 300218 442826 300454
rect 443062 300218 443146 300454
rect 443382 300218 443414 300454
rect 442794 300134 443414 300218
rect 442794 299898 442826 300134
rect 443062 299898 443146 300134
rect 443382 299898 443414 300134
rect 442794 264454 443414 299898
rect 442794 264218 442826 264454
rect 443062 264218 443146 264454
rect 443382 264218 443414 264454
rect 442794 264134 443414 264218
rect 442794 263898 442826 264134
rect 443062 263898 443146 264134
rect 443382 263898 443414 264134
rect 442794 228454 443414 263898
rect 442794 228218 442826 228454
rect 443062 228218 443146 228454
rect 443382 228218 443414 228454
rect 442794 228134 443414 228218
rect 442794 227898 442826 228134
rect 443062 227898 443146 228134
rect 443382 227898 443414 228134
rect 442794 192454 443414 227898
rect 442794 192218 442826 192454
rect 443062 192218 443146 192454
rect 443382 192218 443414 192454
rect 442794 192134 443414 192218
rect 442794 191898 442826 192134
rect 443062 191898 443146 192134
rect 443382 191898 443414 192134
rect 442794 156454 443414 191898
rect 442794 156218 442826 156454
rect 443062 156218 443146 156454
rect 443382 156218 443414 156454
rect 442794 156134 443414 156218
rect 442794 155898 442826 156134
rect 443062 155898 443146 156134
rect 443382 155898 443414 156134
rect 442794 120454 443414 155898
rect 442794 120218 442826 120454
rect 443062 120218 443146 120454
rect 443382 120218 443414 120454
rect 442794 120134 443414 120218
rect 442794 119898 442826 120134
rect 443062 119898 443146 120134
rect 443382 119898 443414 120134
rect 442794 84454 443414 119898
rect 442794 84218 442826 84454
rect 443062 84218 443146 84454
rect 443382 84218 443414 84454
rect 442794 84134 443414 84218
rect 442794 83898 442826 84134
rect 443062 83898 443146 84134
rect 443382 83898 443414 84134
rect 442794 48454 443414 83898
rect 442794 48218 442826 48454
rect 443062 48218 443146 48454
rect 443382 48218 443414 48454
rect 442794 48134 443414 48218
rect 442794 47898 442826 48134
rect 443062 47898 443146 48134
rect 443382 47898 443414 48134
rect 442794 12454 443414 47898
rect 442794 12218 442826 12454
rect 443062 12218 443146 12454
rect 443382 12218 443414 12454
rect 442794 12134 443414 12218
rect 442794 11898 442826 12134
rect 443062 11898 443146 12134
rect 443382 11898 443414 12134
rect 442794 -2266 443414 11898
rect 442794 -2502 442826 -2266
rect 443062 -2502 443146 -2266
rect 443382 -2502 443414 -2266
rect 442794 -2586 443414 -2502
rect 442794 -2822 442826 -2586
rect 443062 -2822 443146 -2586
rect 443382 -2822 443414 -2586
rect 442794 -7654 443414 -2822
rect 447294 484954 447914 498000
rect 447294 484718 447326 484954
rect 447562 484718 447646 484954
rect 447882 484718 447914 484954
rect 447294 484634 447914 484718
rect 447294 484398 447326 484634
rect 447562 484398 447646 484634
rect 447882 484398 447914 484634
rect 447294 448954 447914 484398
rect 447294 448718 447326 448954
rect 447562 448718 447646 448954
rect 447882 448718 447914 448954
rect 447294 448634 447914 448718
rect 447294 448398 447326 448634
rect 447562 448398 447646 448634
rect 447882 448398 447914 448634
rect 447294 412954 447914 448398
rect 447294 412718 447326 412954
rect 447562 412718 447646 412954
rect 447882 412718 447914 412954
rect 447294 412634 447914 412718
rect 447294 412398 447326 412634
rect 447562 412398 447646 412634
rect 447882 412398 447914 412634
rect 447294 376954 447914 412398
rect 447294 376718 447326 376954
rect 447562 376718 447646 376954
rect 447882 376718 447914 376954
rect 447294 376634 447914 376718
rect 447294 376398 447326 376634
rect 447562 376398 447646 376634
rect 447882 376398 447914 376634
rect 447294 340954 447914 376398
rect 447294 340718 447326 340954
rect 447562 340718 447646 340954
rect 447882 340718 447914 340954
rect 447294 340634 447914 340718
rect 447294 340398 447326 340634
rect 447562 340398 447646 340634
rect 447882 340398 447914 340634
rect 447294 304954 447914 340398
rect 447294 304718 447326 304954
rect 447562 304718 447646 304954
rect 447882 304718 447914 304954
rect 447294 304634 447914 304718
rect 447294 304398 447326 304634
rect 447562 304398 447646 304634
rect 447882 304398 447914 304634
rect 447294 268954 447914 304398
rect 447294 268718 447326 268954
rect 447562 268718 447646 268954
rect 447882 268718 447914 268954
rect 447294 268634 447914 268718
rect 447294 268398 447326 268634
rect 447562 268398 447646 268634
rect 447882 268398 447914 268634
rect 447294 232954 447914 268398
rect 447294 232718 447326 232954
rect 447562 232718 447646 232954
rect 447882 232718 447914 232954
rect 447294 232634 447914 232718
rect 447294 232398 447326 232634
rect 447562 232398 447646 232634
rect 447882 232398 447914 232634
rect 447294 196954 447914 232398
rect 447294 196718 447326 196954
rect 447562 196718 447646 196954
rect 447882 196718 447914 196954
rect 447294 196634 447914 196718
rect 447294 196398 447326 196634
rect 447562 196398 447646 196634
rect 447882 196398 447914 196634
rect 447294 160954 447914 196398
rect 447294 160718 447326 160954
rect 447562 160718 447646 160954
rect 447882 160718 447914 160954
rect 447294 160634 447914 160718
rect 447294 160398 447326 160634
rect 447562 160398 447646 160634
rect 447882 160398 447914 160634
rect 447294 124954 447914 160398
rect 447294 124718 447326 124954
rect 447562 124718 447646 124954
rect 447882 124718 447914 124954
rect 447294 124634 447914 124718
rect 447294 124398 447326 124634
rect 447562 124398 447646 124634
rect 447882 124398 447914 124634
rect 447294 88954 447914 124398
rect 447294 88718 447326 88954
rect 447562 88718 447646 88954
rect 447882 88718 447914 88954
rect 447294 88634 447914 88718
rect 447294 88398 447326 88634
rect 447562 88398 447646 88634
rect 447882 88398 447914 88634
rect 447294 52954 447914 88398
rect 447294 52718 447326 52954
rect 447562 52718 447646 52954
rect 447882 52718 447914 52954
rect 447294 52634 447914 52718
rect 447294 52398 447326 52634
rect 447562 52398 447646 52634
rect 447882 52398 447914 52634
rect 447294 16954 447914 52398
rect 447294 16718 447326 16954
rect 447562 16718 447646 16954
rect 447882 16718 447914 16954
rect 447294 16634 447914 16718
rect 447294 16398 447326 16634
rect 447562 16398 447646 16634
rect 447882 16398 447914 16634
rect 447294 -3226 447914 16398
rect 447294 -3462 447326 -3226
rect 447562 -3462 447646 -3226
rect 447882 -3462 447914 -3226
rect 447294 -3546 447914 -3462
rect 447294 -3782 447326 -3546
rect 447562 -3782 447646 -3546
rect 447882 -3782 447914 -3546
rect 447294 -7654 447914 -3782
rect 451794 489454 452414 498000
rect 451794 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 452414 489454
rect 451794 489134 452414 489218
rect 451794 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 452414 489134
rect 451794 453454 452414 488898
rect 451794 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 452414 453454
rect 451794 453134 452414 453218
rect 451794 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 452414 453134
rect 451794 417454 452414 452898
rect 451794 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 452414 417454
rect 451794 417134 452414 417218
rect 451794 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 452414 417134
rect 451794 381454 452414 416898
rect 451794 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 452414 381454
rect 451794 381134 452414 381218
rect 451794 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 452414 381134
rect 451794 345454 452414 380898
rect 451794 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 452414 345454
rect 451794 345134 452414 345218
rect 451794 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 452414 345134
rect 451794 309454 452414 344898
rect 451794 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 452414 309454
rect 451794 309134 452414 309218
rect 451794 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 452414 309134
rect 451794 273454 452414 308898
rect 451794 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 452414 273454
rect 451794 273134 452414 273218
rect 451794 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 452414 273134
rect 451794 237454 452414 272898
rect 451794 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 452414 237454
rect 451794 237134 452414 237218
rect 451794 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 452414 237134
rect 451794 201454 452414 236898
rect 451794 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 452414 201454
rect 451794 201134 452414 201218
rect 451794 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 452414 201134
rect 451794 165454 452414 200898
rect 451794 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 452414 165454
rect 451794 165134 452414 165218
rect 451794 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 452414 165134
rect 451794 129454 452414 164898
rect 451794 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 452414 129454
rect 451794 129134 452414 129218
rect 451794 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 452414 129134
rect 451794 93454 452414 128898
rect 451794 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 452414 93454
rect 451794 93134 452414 93218
rect 451794 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 452414 93134
rect 451794 57454 452414 92898
rect 451794 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 452414 57454
rect 451794 57134 452414 57218
rect 451794 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 452414 57134
rect 451794 21454 452414 56898
rect 451794 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 452414 21454
rect 451794 21134 452414 21218
rect 451794 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 452414 21134
rect 451794 -4186 452414 20898
rect 451794 -4422 451826 -4186
rect 452062 -4422 452146 -4186
rect 452382 -4422 452414 -4186
rect 451794 -4506 452414 -4422
rect 451794 -4742 451826 -4506
rect 452062 -4742 452146 -4506
rect 452382 -4742 452414 -4506
rect 451794 -7654 452414 -4742
rect 456294 493954 456914 498000
rect 456294 493718 456326 493954
rect 456562 493718 456646 493954
rect 456882 493718 456914 493954
rect 456294 493634 456914 493718
rect 456294 493398 456326 493634
rect 456562 493398 456646 493634
rect 456882 493398 456914 493634
rect 456294 457954 456914 493398
rect 456294 457718 456326 457954
rect 456562 457718 456646 457954
rect 456882 457718 456914 457954
rect 456294 457634 456914 457718
rect 456294 457398 456326 457634
rect 456562 457398 456646 457634
rect 456882 457398 456914 457634
rect 456294 421954 456914 457398
rect 456294 421718 456326 421954
rect 456562 421718 456646 421954
rect 456882 421718 456914 421954
rect 456294 421634 456914 421718
rect 456294 421398 456326 421634
rect 456562 421398 456646 421634
rect 456882 421398 456914 421634
rect 456294 385954 456914 421398
rect 456294 385718 456326 385954
rect 456562 385718 456646 385954
rect 456882 385718 456914 385954
rect 456294 385634 456914 385718
rect 456294 385398 456326 385634
rect 456562 385398 456646 385634
rect 456882 385398 456914 385634
rect 456294 349954 456914 385398
rect 456294 349718 456326 349954
rect 456562 349718 456646 349954
rect 456882 349718 456914 349954
rect 456294 349634 456914 349718
rect 456294 349398 456326 349634
rect 456562 349398 456646 349634
rect 456882 349398 456914 349634
rect 456294 313954 456914 349398
rect 456294 313718 456326 313954
rect 456562 313718 456646 313954
rect 456882 313718 456914 313954
rect 456294 313634 456914 313718
rect 456294 313398 456326 313634
rect 456562 313398 456646 313634
rect 456882 313398 456914 313634
rect 456294 277954 456914 313398
rect 456294 277718 456326 277954
rect 456562 277718 456646 277954
rect 456882 277718 456914 277954
rect 456294 277634 456914 277718
rect 456294 277398 456326 277634
rect 456562 277398 456646 277634
rect 456882 277398 456914 277634
rect 456294 241954 456914 277398
rect 456294 241718 456326 241954
rect 456562 241718 456646 241954
rect 456882 241718 456914 241954
rect 456294 241634 456914 241718
rect 456294 241398 456326 241634
rect 456562 241398 456646 241634
rect 456882 241398 456914 241634
rect 456294 205954 456914 241398
rect 456294 205718 456326 205954
rect 456562 205718 456646 205954
rect 456882 205718 456914 205954
rect 456294 205634 456914 205718
rect 456294 205398 456326 205634
rect 456562 205398 456646 205634
rect 456882 205398 456914 205634
rect 456294 169954 456914 205398
rect 456294 169718 456326 169954
rect 456562 169718 456646 169954
rect 456882 169718 456914 169954
rect 456294 169634 456914 169718
rect 456294 169398 456326 169634
rect 456562 169398 456646 169634
rect 456882 169398 456914 169634
rect 456294 133954 456914 169398
rect 456294 133718 456326 133954
rect 456562 133718 456646 133954
rect 456882 133718 456914 133954
rect 456294 133634 456914 133718
rect 456294 133398 456326 133634
rect 456562 133398 456646 133634
rect 456882 133398 456914 133634
rect 456294 97954 456914 133398
rect 456294 97718 456326 97954
rect 456562 97718 456646 97954
rect 456882 97718 456914 97954
rect 456294 97634 456914 97718
rect 456294 97398 456326 97634
rect 456562 97398 456646 97634
rect 456882 97398 456914 97634
rect 456294 61954 456914 97398
rect 456294 61718 456326 61954
rect 456562 61718 456646 61954
rect 456882 61718 456914 61954
rect 456294 61634 456914 61718
rect 456294 61398 456326 61634
rect 456562 61398 456646 61634
rect 456882 61398 456914 61634
rect 456294 25954 456914 61398
rect 456294 25718 456326 25954
rect 456562 25718 456646 25954
rect 456882 25718 456914 25954
rect 456294 25634 456914 25718
rect 456294 25398 456326 25634
rect 456562 25398 456646 25634
rect 456882 25398 456914 25634
rect 456294 -5146 456914 25398
rect 456294 -5382 456326 -5146
rect 456562 -5382 456646 -5146
rect 456882 -5382 456914 -5146
rect 456294 -5466 456914 -5382
rect 456294 -5702 456326 -5466
rect 456562 -5702 456646 -5466
rect 456882 -5702 456914 -5466
rect 456294 -7654 456914 -5702
rect 460794 462454 461414 498000
rect 460794 462218 460826 462454
rect 461062 462218 461146 462454
rect 461382 462218 461414 462454
rect 460794 462134 461414 462218
rect 460794 461898 460826 462134
rect 461062 461898 461146 462134
rect 461382 461898 461414 462134
rect 460794 426454 461414 461898
rect 460794 426218 460826 426454
rect 461062 426218 461146 426454
rect 461382 426218 461414 426454
rect 460794 426134 461414 426218
rect 460794 425898 460826 426134
rect 461062 425898 461146 426134
rect 461382 425898 461414 426134
rect 460794 390454 461414 425898
rect 460794 390218 460826 390454
rect 461062 390218 461146 390454
rect 461382 390218 461414 390454
rect 460794 390134 461414 390218
rect 460794 389898 460826 390134
rect 461062 389898 461146 390134
rect 461382 389898 461414 390134
rect 460794 354454 461414 389898
rect 460794 354218 460826 354454
rect 461062 354218 461146 354454
rect 461382 354218 461414 354454
rect 460794 354134 461414 354218
rect 460794 353898 460826 354134
rect 461062 353898 461146 354134
rect 461382 353898 461414 354134
rect 460794 318454 461414 353898
rect 460794 318218 460826 318454
rect 461062 318218 461146 318454
rect 461382 318218 461414 318454
rect 460794 318134 461414 318218
rect 460794 317898 460826 318134
rect 461062 317898 461146 318134
rect 461382 317898 461414 318134
rect 460794 282454 461414 317898
rect 460794 282218 460826 282454
rect 461062 282218 461146 282454
rect 461382 282218 461414 282454
rect 460794 282134 461414 282218
rect 460794 281898 460826 282134
rect 461062 281898 461146 282134
rect 461382 281898 461414 282134
rect 460794 246454 461414 281898
rect 460794 246218 460826 246454
rect 461062 246218 461146 246454
rect 461382 246218 461414 246454
rect 460794 246134 461414 246218
rect 460794 245898 460826 246134
rect 461062 245898 461146 246134
rect 461382 245898 461414 246134
rect 460794 210454 461414 245898
rect 460794 210218 460826 210454
rect 461062 210218 461146 210454
rect 461382 210218 461414 210454
rect 460794 210134 461414 210218
rect 460794 209898 460826 210134
rect 461062 209898 461146 210134
rect 461382 209898 461414 210134
rect 460794 174454 461414 209898
rect 460794 174218 460826 174454
rect 461062 174218 461146 174454
rect 461382 174218 461414 174454
rect 460794 174134 461414 174218
rect 460794 173898 460826 174134
rect 461062 173898 461146 174134
rect 461382 173898 461414 174134
rect 460794 138454 461414 173898
rect 460794 138218 460826 138454
rect 461062 138218 461146 138454
rect 461382 138218 461414 138454
rect 460794 138134 461414 138218
rect 460794 137898 460826 138134
rect 461062 137898 461146 138134
rect 461382 137898 461414 138134
rect 460794 102454 461414 137898
rect 460794 102218 460826 102454
rect 461062 102218 461146 102454
rect 461382 102218 461414 102454
rect 460794 102134 461414 102218
rect 460794 101898 460826 102134
rect 461062 101898 461146 102134
rect 461382 101898 461414 102134
rect 460794 66454 461414 101898
rect 460794 66218 460826 66454
rect 461062 66218 461146 66454
rect 461382 66218 461414 66454
rect 460794 66134 461414 66218
rect 460794 65898 460826 66134
rect 461062 65898 461146 66134
rect 461382 65898 461414 66134
rect 460794 30454 461414 65898
rect 460794 30218 460826 30454
rect 461062 30218 461146 30454
rect 461382 30218 461414 30454
rect 460794 30134 461414 30218
rect 460794 29898 460826 30134
rect 461062 29898 461146 30134
rect 461382 29898 461414 30134
rect 460794 -6106 461414 29898
rect 460794 -6342 460826 -6106
rect 461062 -6342 461146 -6106
rect 461382 -6342 461414 -6106
rect 460794 -6426 461414 -6342
rect 460794 -6662 460826 -6426
rect 461062 -6662 461146 -6426
rect 461382 -6662 461414 -6426
rect 460794 -7654 461414 -6662
rect 465294 466954 465914 498000
rect 465294 466718 465326 466954
rect 465562 466718 465646 466954
rect 465882 466718 465914 466954
rect 465294 466634 465914 466718
rect 465294 466398 465326 466634
rect 465562 466398 465646 466634
rect 465882 466398 465914 466634
rect 465294 430954 465914 466398
rect 465294 430718 465326 430954
rect 465562 430718 465646 430954
rect 465882 430718 465914 430954
rect 465294 430634 465914 430718
rect 465294 430398 465326 430634
rect 465562 430398 465646 430634
rect 465882 430398 465914 430634
rect 465294 394954 465914 430398
rect 465294 394718 465326 394954
rect 465562 394718 465646 394954
rect 465882 394718 465914 394954
rect 465294 394634 465914 394718
rect 465294 394398 465326 394634
rect 465562 394398 465646 394634
rect 465882 394398 465914 394634
rect 465294 358954 465914 394398
rect 465294 358718 465326 358954
rect 465562 358718 465646 358954
rect 465882 358718 465914 358954
rect 465294 358634 465914 358718
rect 465294 358398 465326 358634
rect 465562 358398 465646 358634
rect 465882 358398 465914 358634
rect 465294 322954 465914 358398
rect 465294 322718 465326 322954
rect 465562 322718 465646 322954
rect 465882 322718 465914 322954
rect 465294 322634 465914 322718
rect 465294 322398 465326 322634
rect 465562 322398 465646 322634
rect 465882 322398 465914 322634
rect 465294 286954 465914 322398
rect 465294 286718 465326 286954
rect 465562 286718 465646 286954
rect 465882 286718 465914 286954
rect 465294 286634 465914 286718
rect 465294 286398 465326 286634
rect 465562 286398 465646 286634
rect 465882 286398 465914 286634
rect 465294 250954 465914 286398
rect 465294 250718 465326 250954
rect 465562 250718 465646 250954
rect 465882 250718 465914 250954
rect 465294 250634 465914 250718
rect 465294 250398 465326 250634
rect 465562 250398 465646 250634
rect 465882 250398 465914 250634
rect 465294 214954 465914 250398
rect 465294 214718 465326 214954
rect 465562 214718 465646 214954
rect 465882 214718 465914 214954
rect 465294 214634 465914 214718
rect 465294 214398 465326 214634
rect 465562 214398 465646 214634
rect 465882 214398 465914 214634
rect 465294 178954 465914 214398
rect 465294 178718 465326 178954
rect 465562 178718 465646 178954
rect 465882 178718 465914 178954
rect 465294 178634 465914 178718
rect 465294 178398 465326 178634
rect 465562 178398 465646 178634
rect 465882 178398 465914 178634
rect 465294 142954 465914 178398
rect 465294 142718 465326 142954
rect 465562 142718 465646 142954
rect 465882 142718 465914 142954
rect 465294 142634 465914 142718
rect 465294 142398 465326 142634
rect 465562 142398 465646 142634
rect 465882 142398 465914 142634
rect 465294 106954 465914 142398
rect 465294 106718 465326 106954
rect 465562 106718 465646 106954
rect 465882 106718 465914 106954
rect 465294 106634 465914 106718
rect 465294 106398 465326 106634
rect 465562 106398 465646 106634
rect 465882 106398 465914 106634
rect 465294 70954 465914 106398
rect 465294 70718 465326 70954
rect 465562 70718 465646 70954
rect 465882 70718 465914 70954
rect 465294 70634 465914 70718
rect 465294 70398 465326 70634
rect 465562 70398 465646 70634
rect 465882 70398 465914 70634
rect 465294 34954 465914 70398
rect 465294 34718 465326 34954
rect 465562 34718 465646 34954
rect 465882 34718 465914 34954
rect 465294 34634 465914 34718
rect 465294 34398 465326 34634
rect 465562 34398 465646 34634
rect 465882 34398 465914 34634
rect 465294 -7066 465914 34398
rect 465294 -7302 465326 -7066
rect 465562 -7302 465646 -7066
rect 465882 -7302 465914 -7066
rect 465294 -7386 465914 -7302
rect 465294 -7622 465326 -7386
rect 465562 -7622 465646 -7386
rect 465882 -7622 465914 -7386
rect 465294 -7654 465914 -7622
rect 469794 471454 470414 498000
rect 469794 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 470414 471454
rect 469794 471134 470414 471218
rect 469794 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 470414 471134
rect 469794 435454 470414 470898
rect 469794 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 470414 435454
rect 469794 435134 470414 435218
rect 469794 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 470414 435134
rect 469794 399454 470414 434898
rect 469794 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 470414 399454
rect 469794 399134 470414 399218
rect 469794 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 470414 399134
rect 469794 363454 470414 398898
rect 469794 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 470414 363454
rect 469794 363134 470414 363218
rect 469794 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 470414 363134
rect 469794 327454 470414 362898
rect 469794 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 470414 327454
rect 469794 327134 470414 327218
rect 469794 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 470414 327134
rect 469794 291454 470414 326898
rect 469794 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 470414 291454
rect 469794 291134 470414 291218
rect 469794 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 470414 291134
rect 469794 255454 470414 290898
rect 469794 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 470414 255454
rect 469794 255134 470414 255218
rect 469794 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 470414 255134
rect 469794 219454 470414 254898
rect 469794 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 470414 219454
rect 469794 219134 470414 219218
rect 469794 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 470414 219134
rect 469794 183454 470414 218898
rect 469794 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 470414 183454
rect 469794 183134 470414 183218
rect 469794 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 470414 183134
rect 469794 147454 470414 182898
rect 469794 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 470414 147454
rect 469794 147134 470414 147218
rect 469794 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 470414 147134
rect 469794 111454 470414 146898
rect 469794 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 470414 111454
rect 469794 111134 470414 111218
rect 469794 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 470414 111134
rect 469794 75454 470414 110898
rect 469794 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 470414 75454
rect 469794 75134 470414 75218
rect 469794 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 470414 75134
rect 469794 39454 470414 74898
rect 469794 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 470414 39454
rect 469794 39134 470414 39218
rect 469794 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 470414 39134
rect 469794 3454 470414 38898
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -7654 470414 -902
rect 474294 475954 474914 511398
rect 474294 475718 474326 475954
rect 474562 475718 474646 475954
rect 474882 475718 474914 475954
rect 474294 475634 474914 475718
rect 474294 475398 474326 475634
rect 474562 475398 474646 475634
rect 474882 475398 474914 475634
rect 474294 439954 474914 475398
rect 474294 439718 474326 439954
rect 474562 439718 474646 439954
rect 474882 439718 474914 439954
rect 474294 439634 474914 439718
rect 474294 439398 474326 439634
rect 474562 439398 474646 439634
rect 474882 439398 474914 439634
rect 474294 403954 474914 439398
rect 474294 403718 474326 403954
rect 474562 403718 474646 403954
rect 474882 403718 474914 403954
rect 474294 403634 474914 403718
rect 474294 403398 474326 403634
rect 474562 403398 474646 403634
rect 474882 403398 474914 403634
rect 474294 367954 474914 403398
rect 474294 367718 474326 367954
rect 474562 367718 474646 367954
rect 474882 367718 474914 367954
rect 474294 367634 474914 367718
rect 474294 367398 474326 367634
rect 474562 367398 474646 367634
rect 474882 367398 474914 367634
rect 474294 331954 474914 367398
rect 474294 331718 474326 331954
rect 474562 331718 474646 331954
rect 474882 331718 474914 331954
rect 474294 331634 474914 331718
rect 474294 331398 474326 331634
rect 474562 331398 474646 331634
rect 474882 331398 474914 331634
rect 474294 295954 474914 331398
rect 474294 295718 474326 295954
rect 474562 295718 474646 295954
rect 474882 295718 474914 295954
rect 474294 295634 474914 295718
rect 474294 295398 474326 295634
rect 474562 295398 474646 295634
rect 474882 295398 474914 295634
rect 474294 259954 474914 295398
rect 474294 259718 474326 259954
rect 474562 259718 474646 259954
rect 474882 259718 474914 259954
rect 474294 259634 474914 259718
rect 474294 259398 474326 259634
rect 474562 259398 474646 259634
rect 474882 259398 474914 259634
rect 474294 223954 474914 259398
rect 474294 223718 474326 223954
rect 474562 223718 474646 223954
rect 474882 223718 474914 223954
rect 474294 223634 474914 223718
rect 474294 223398 474326 223634
rect 474562 223398 474646 223634
rect 474882 223398 474914 223634
rect 474294 187954 474914 223398
rect 474294 187718 474326 187954
rect 474562 187718 474646 187954
rect 474882 187718 474914 187954
rect 474294 187634 474914 187718
rect 474294 187398 474326 187634
rect 474562 187398 474646 187634
rect 474882 187398 474914 187634
rect 474294 151954 474914 187398
rect 474294 151718 474326 151954
rect 474562 151718 474646 151954
rect 474882 151718 474914 151954
rect 474294 151634 474914 151718
rect 474294 151398 474326 151634
rect 474562 151398 474646 151634
rect 474882 151398 474914 151634
rect 474294 115954 474914 151398
rect 474294 115718 474326 115954
rect 474562 115718 474646 115954
rect 474882 115718 474914 115954
rect 474294 115634 474914 115718
rect 474294 115398 474326 115634
rect 474562 115398 474646 115634
rect 474882 115398 474914 115634
rect 474294 79954 474914 115398
rect 474294 79718 474326 79954
rect 474562 79718 474646 79954
rect 474882 79718 474914 79954
rect 474294 79634 474914 79718
rect 474294 79398 474326 79634
rect 474562 79398 474646 79634
rect 474882 79398 474914 79634
rect 474294 43954 474914 79398
rect 474294 43718 474326 43954
rect 474562 43718 474646 43954
rect 474882 43718 474914 43954
rect 474294 43634 474914 43718
rect 474294 43398 474326 43634
rect 474562 43398 474646 43634
rect 474882 43398 474914 43634
rect 474294 7954 474914 43398
rect 474294 7718 474326 7954
rect 474562 7718 474646 7954
rect 474882 7718 474914 7954
rect 474294 7634 474914 7718
rect 474294 7398 474326 7634
rect 474562 7398 474646 7634
rect 474882 7398 474914 7634
rect 474294 -1306 474914 7398
rect 474294 -1542 474326 -1306
rect 474562 -1542 474646 -1306
rect 474882 -1542 474914 -1306
rect 474294 -1626 474914 -1542
rect 474294 -1862 474326 -1626
rect 474562 -1862 474646 -1626
rect 474882 -1862 474914 -1626
rect 474294 -7654 474914 -1862
rect 478794 706758 479414 711590
rect 478794 706522 478826 706758
rect 479062 706522 479146 706758
rect 479382 706522 479414 706758
rect 478794 706438 479414 706522
rect 478794 706202 478826 706438
rect 479062 706202 479146 706438
rect 479382 706202 479414 706438
rect 478794 696454 479414 706202
rect 478794 696218 478826 696454
rect 479062 696218 479146 696454
rect 479382 696218 479414 696454
rect 478794 696134 479414 696218
rect 478794 695898 478826 696134
rect 479062 695898 479146 696134
rect 479382 695898 479414 696134
rect 478794 660454 479414 695898
rect 478794 660218 478826 660454
rect 479062 660218 479146 660454
rect 479382 660218 479414 660454
rect 478794 660134 479414 660218
rect 478794 659898 478826 660134
rect 479062 659898 479146 660134
rect 479382 659898 479414 660134
rect 478794 624454 479414 659898
rect 478794 624218 478826 624454
rect 479062 624218 479146 624454
rect 479382 624218 479414 624454
rect 478794 624134 479414 624218
rect 478794 623898 478826 624134
rect 479062 623898 479146 624134
rect 479382 623898 479414 624134
rect 478794 588454 479414 623898
rect 478794 588218 478826 588454
rect 479062 588218 479146 588454
rect 479382 588218 479414 588454
rect 478794 588134 479414 588218
rect 478794 587898 478826 588134
rect 479062 587898 479146 588134
rect 479382 587898 479414 588134
rect 478794 552454 479414 587898
rect 478794 552218 478826 552454
rect 479062 552218 479146 552454
rect 479382 552218 479414 552454
rect 478794 552134 479414 552218
rect 478794 551898 478826 552134
rect 479062 551898 479146 552134
rect 479382 551898 479414 552134
rect 478794 516454 479414 551898
rect 478794 516218 478826 516454
rect 479062 516218 479146 516454
rect 479382 516218 479414 516454
rect 478794 516134 479414 516218
rect 478794 515898 478826 516134
rect 479062 515898 479146 516134
rect 479382 515898 479414 516134
rect 478794 480454 479414 515898
rect 478794 480218 478826 480454
rect 479062 480218 479146 480454
rect 479382 480218 479414 480454
rect 478794 480134 479414 480218
rect 478794 479898 478826 480134
rect 479062 479898 479146 480134
rect 479382 479898 479414 480134
rect 478794 444454 479414 479898
rect 478794 444218 478826 444454
rect 479062 444218 479146 444454
rect 479382 444218 479414 444454
rect 478794 444134 479414 444218
rect 478794 443898 478826 444134
rect 479062 443898 479146 444134
rect 479382 443898 479414 444134
rect 478794 408454 479414 443898
rect 478794 408218 478826 408454
rect 479062 408218 479146 408454
rect 479382 408218 479414 408454
rect 478794 408134 479414 408218
rect 478794 407898 478826 408134
rect 479062 407898 479146 408134
rect 479382 407898 479414 408134
rect 478794 372454 479414 407898
rect 478794 372218 478826 372454
rect 479062 372218 479146 372454
rect 479382 372218 479414 372454
rect 478794 372134 479414 372218
rect 478794 371898 478826 372134
rect 479062 371898 479146 372134
rect 479382 371898 479414 372134
rect 478794 336454 479414 371898
rect 478794 336218 478826 336454
rect 479062 336218 479146 336454
rect 479382 336218 479414 336454
rect 478794 336134 479414 336218
rect 478794 335898 478826 336134
rect 479062 335898 479146 336134
rect 479382 335898 479414 336134
rect 478794 300454 479414 335898
rect 478794 300218 478826 300454
rect 479062 300218 479146 300454
rect 479382 300218 479414 300454
rect 478794 300134 479414 300218
rect 478794 299898 478826 300134
rect 479062 299898 479146 300134
rect 479382 299898 479414 300134
rect 478794 264454 479414 299898
rect 478794 264218 478826 264454
rect 479062 264218 479146 264454
rect 479382 264218 479414 264454
rect 478794 264134 479414 264218
rect 478794 263898 478826 264134
rect 479062 263898 479146 264134
rect 479382 263898 479414 264134
rect 478794 228454 479414 263898
rect 478794 228218 478826 228454
rect 479062 228218 479146 228454
rect 479382 228218 479414 228454
rect 478794 228134 479414 228218
rect 478794 227898 478826 228134
rect 479062 227898 479146 228134
rect 479382 227898 479414 228134
rect 478794 192454 479414 227898
rect 478794 192218 478826 192454
rect 479062 192218 479146 192454
rect 479382 192218 479414 192454
rect 478794 192134 479414 192218
rect 478794 191898 478826 192134
rect 479062 191898 479146 192134
rect 479382 191898 479414 192134
rect 478794 156454 479414 191898
rect 478794 156218 478826 156454
rect 479062 156218 479146 156454
rect 479382 156218 479414 156454
rect 478794 156134 479414 156218
rect 478794 155898 478826 156134
rect 479062 155898 479146 156134
rect 479382 155898 479414 156134
rect 478794 120454 479414 155898
rect 478794 120218 478826 120454
rect 479062 120218 479146 120454
rect 479382 120218 479414 120454
rect 478794 120134 479414 120218
rect 478794 119898 478826 120134
rect 479062 119898 479146 120134
rect 479382 119898 479414 120134
rect 478794 84454 479414 119898
rect 478794 84218 478826 84454
rect 479062 84218 479146 84454
rect 479382 84218 479414 84454
rect 478794 84134 479414 84218
rect 478794 83898 478826 84134
rect 479062 83898 479146 84134
rect 479382 83898 479414 84134
rect 478794 48454 479414 83898
rect 478794 48218 478826 48454
rect 479062 48218 479146 48454
rect 479382 48218 479414 48454
rect 478794 48134 479414 48218
rect 478794 47898 478826 48134
rect 479062 47898 479146 48134
rect 479382 47898 479414 48134
rect 478794 12454 479414 47898
rect 478794 12218 478826 12454
rect 479062 12218 479146 12454
rect 479382 12218 479414 12454
rect 478794 12134 479414 12218
rect 478794 11898 478826 12134
rect 479062 11898 479146 12134
rect 479382 11898 479414 12134
rect 478794 -2266 479414 11898
rect 478794 -2502 478826 -2266
rect 479062 -2502 479146 -2266
rect 479382 -2502 479414 -2266
rect 478794 -2586 479414 -2502
rect 478794 -2822 478826 -2586
rect 479062 -2822 479146 -2586
rect 479382 -2822 479414 -2586
rect 478794 -7654 479414 -2822
rect 483294 707718 483914 711590
rect 483294 707482 483326 707718
rect 483562 707482 483646 707718
rect 483882 707482 483914 707718
rect 483294 707398 483914 707482
rect 483294 707162 483326 707398
rect 483562 707162 483646 707398
rect 483882 707162 483914 707398
rect 483294 700954 483914 707162
rect 483294 700718 483326 700954
rect 483562 700718 483646 700954
rect 483882 700718 483914 700954
rect 483294 700634 483914 700718
rect 483294 700398 483326 700634
rect 483562 700398 483646 700634
rect 483882 700398 483914 700634
rect 483294 664954 483914 700398
rect 483294 664718 483326 664954
rect 483562 664718 483646 664954
rect 483882 664718 483914 664954
rect 483294 664634 483914 664718
rect 483294 664398 483326 664634
rect 483562 664398 483646 664634
rect 483882 664398 483914 664634
rect 483294 628954 483914 664398
rect 483294 628718 483326 628954
rect 483562 628718 483646 628954
rect 483882 628718 483914 628954
rect 483294 628634 483914 628718
rect 483294 628398 483326 628634
rect 483562 628398 483646 628634
rect 483882 628398 483914 628634
rect 483294 592954 483914 628398
rect 483294 592718 483326 592954
rect 483562 592718 483646 592954
rect 483882 592718 483914 592954
rect 483294 592634 483914 592718
rect 483294 592398 483326 592634
rect 483562 592398 483646 592634
rect 483882 592398 483914 592634
rect 483294 556954 483914 592398
rect 483294 556718 483326 556954
rect 483562 556718 483646 556954
rect 483882 556718 483914 556954
rect 483294 556634 483914 556718
rect 483294 556398 483326 556634
rect 483562 556398 483646 556634
rect 483882 556398 483914 556634
rect 483294 520954 483914 556398
rect 483294 520718 483326 520954
rect 483562 520718 483646 520954
rect 483882 520718 483914 520954
rect 483294 520634 483914 520718
rect 483294 520398 483326 520634
rect 483562 520398 483646 520634
rect 483882 520398 483914 520634
rect 483294 484954 483914 520398
rect 483294 484718 483326 484954
rect 483562 484718 483646 484954
rect 483882 484718 483914 484954
rect 483294 484634 483914 484718
rect 483294 484398 483326 484634
rect 483562 484398 483646 484634
rect 483882 484398 483914 484634
rect 483294 448954 483914 484398
rect 483294 448718 483326 448954
rect 483562 448718 483646 448954
rect 483882 448718 483914 448954
rect 483294 448634 483914 448718
rect 483294 448398 483326 448634
rect 483562 448398 483646 448634
rect 483882 448398 483914 448634
rect 483294 412954 483914 448398
rect 483294 412718 483326 412954
rect 483562 412718 483646 412954
rect 483882 412718 483914 412954
rect 483294 412634 483914 412718
rect 483294 412398 483326 412634
rect 483562 412398 483646 412634
rect 483882 412398 483914 412634
rect 483294 376954 483914 412398
rect 483294 376718 483326 376954
rect 483562 376718 483646 376954
rect 483882 376718 483914 376954
rect 483294 376634 483914 376718
rect 483294 376398 483326 376634
rect 483562 376398 483646 376634
rect 483882 376398 483914 376634
rect 483294 340954 483914 376398
rect 483294 340718 483326 340954
rect 483562 340718 483646 340954
rect 483882 340718 483914 340954
rect 483294 340634 483914 340718
rect 483294 340398 483326 340634
rect 483562 340398 483646 340634
rect 483882 340398 483914 340634
rect 483294 304954 483914 340398
rect 483294 304718 483326 304954
rect 483562 304718 483646 304954
rect 483882 304718 483914 304954
rect 483294 304634 483914 304718
rect 483294 304398 483326 304634
rect 483562 304398 483646 304634
rect 483882 304398 483914 304634
rect 483294 268954 483914 304398
rect 483294 268718 483326 268954
rect 483562 268718 483646 268954
rect 483882 268718 483914 268954
rect 483294 268634 483914 268718
rect 483294 268398 483326 268634
rect 483562 268398 483646 268634
rect 483882 268398 483914 268634
rect 483294 232954 483914 268398
rect 483294 232718 483326 232954
rect 483562 232718 483646 232954
rect 483882 232718 483914 232954
rect 483294 232634 483914 232718
rect 483294 232398 483326 232634
rect 483562 232398 483646 232634
rect 483882 232398 483914 232634
rect 483294 196954 483914 232398
rect 483294 196718 483326 196954
rect 483562 196718 483646 196954
rect 483882 196718 483914 196954
rect 483294 196634 483914 196718
rect 483294 196398 483326 196634
rect 483562 196398 483646 196634
rect 483882 196398 483914 196634
rect 483294 160954 483914 196398
rect 483294 160718 483326 160954
rect 483562 160718 483646 160954
rect 483882 160718 483914 160954
rect 483294 160634 483914 160718
rect 483294 160398 483326 160634
rect 483562 160398 483646 160634
rect 483882 160398 483914 160634
rect 483294 124954 483914 160398
rect 483294 124718 483326 124954
rect 483562 124718 483646 124954
rect 483882 124718 483914 124954
rect 483294 124634 483914 124718
rect 483294 124398 483326 124634
rect 483562 124398 483646 124634
rect 483882 124398 483914 124634
rect 483294 88954 483914 124398
rect 483294 88718 483326 88954
rect 483562 88718 483646 88954
rect 483882 88718 483914 88954
rect 483294 88634 483914 88718
rect 483294 88398 483326 88634
rect 483562 88398 483646 88634
rect 483882 88398 483914 88634
rect 483294 52954 483914 88398
rect 483294 52718 483326 52954
rect 483562 52718 483646 52954
rect 483882 52718 483914 52954
rect 483294 52634 483914 52718
rect 483294 52398 483326 52634
rect 483562 52398 483646 52634
rect 483882 52398 483914 52634
rect 483294 16954 483914 52398
rect 483294 16718 483326 16954
rect 483562 16718 483646 16954
rect 483882 16718 483914 16954
rect 483294 16634 483914 16718
rect 483294 16398 483326 16634
rect 483562 16398 483646 16634
rect 483882 16398 483914 16634
rect 483294 -3226 483914 16398
rect 483294 -3462 483326 -3226
rect 483562 -3462 483646 -3226
rect 483882 -3462 483914 -3226
rect 483294 -3546 483914 -3462
rect 483294 -3782 483326 -3546
rect 483562 -3782 483646 -3546
rect 483882 -3782 483914 -3546
rect 483294 -7654 483914 -3782
rect 487794 708678 488414 711590
rect 487794 708442 487826 708678
rect 488062 708442 488146 708678
rect 488382 708442 488414 708678
rect 487794 708358 488414 708442
rect 487794 708122 487826 708358
rect 488062 708122 488146 708358
rect 488382 708122 488414 708358
rect 487794 669454 488414 708122
rect 487794 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 488414 669454
rect 487794 669134 488414 669218
rect 487794 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 488414 669134
rect 487794 633454 488414 668898
rect 487794 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 488414 633454
rect 487794 633134 488414 633218
rect 487794 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 488414 633134
rect 487794 597454 488414 632898
rect 487794 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 488414 597454
rect 487794 597134 488414 597218
rect 487794 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 488414 597134
rect 487794 561454 488414 596898
rect 487794 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 488414 561454
rect 487794 561134 488414 561218
rect 487794 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 488414 561134
rect 487794 525454 488414 560898
rect 487794 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 488414 525454
rect 487794 525134 488414 525218
rect 487794 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 488414 525134
rect 487794 489454 488414 524898
rect 487794 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 488414 489454
rect 487794 489134 488414 489218
rect 487794 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 488414 489134
rect 487794 453454 488414 488898
rect 487794 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 488414 453454
rect 487794 453134 488414 453218
rect 487794 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 488414 453134
rect 487794 417454 488414 452898
rect 487794 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 488414 417454
rect 487794 417134 488414 417218
rect 487794 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 488414 417134
rect 487794 381454 488414 416898
rect 487794 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 488414 381454
rect 487794 381134 488414 381218
rect 487794 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 488414 381134
rect 487794 345454 488414 380898
rect 487794 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 488414 345454
rect 487794 345134 488414 345218
rect 487794 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 488414 345134
rect 487794 309454 488414 344898
rect 487794 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 488414 309454
rect 487794 309134 488414 309218
rect 487794 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 488414 309134
rect 487794 273454 488414 308898
rect 487794 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 488414 273454
rect 487794 273134 488414 273218
rect 487794 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 488414 273134
rect 487794 237454 488414 272898
rect 487794 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 488414 237454
rect 487794 237134 488414 237218
rect 487794 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 488414 237134
rect 487794 201454 488414 236898
rect 487794 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 488414 201454
rect 487794 201134 488414 201218
rect 487794 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 488414 201134
rect 487794 165454 488414 200898
rect 487794 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 488414 165454
rect 487794 165134 488414 165218
rect 487794 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 488414 165134
rect 487794 129454 488414 164898
rect 487794 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 488414 129454
rect 487794 129134 488414 129218
rect 487794 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 488414 129134
rect 487794 93454 488414 128898
rect 487794 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 488414 93454
rect 487794 93134 488414 93218
rect 487794 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 488414 93134
rect 487794 57454 488414 92898
rect 487794 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 488414 57454
rect 487794 57134 488414 57218
rect 487794 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 488414 57134
rect 487794 21454 488414 56898
rect 487794 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 488414 21454
rect 487794 21134 488414 21218
rect 487794 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 488414 21134
rect 487794 -4186 488414 20898
rect 487794 -4422 487826 -4186
rect 488062 -4422 488146 -4186
rect 488382 -4422 488414 -4186
rect 487794 -4506 488414 -4422
rect 487794 -4742 487826 -4506
rect 488062 -4742 488146 -4506
rect 488382 -4742 488414 -4506
rect 487794 -7654 488414 -4742
rect 492294 709638 492914 711590
rect 492294 709402 492326 709638
rect 492562 709402 492646 709638
rect 492882 709402 492914 709638
rect 492294 709318 492914 709402
rect 492294 709082 492326 709318
rect 492562 709082 492646 709318
rect 492882 709082 492914 709318
rect 492294 673954 492914 709082
rect 492294 673718 492326 673954
rect 492562 673718 492646 673954
rect 492882 673718 492914 673954
rect 492294 673634 492914 673718
rect 492294 673398 492326 673634
rect 492562 673398 492646 673634
rect 492882 673398 492914 673634
rect 492294 637954 492914 673398
rect 492294 637718 492326 637954
rect 492562 637718 492646 637954
rect 492882 637718 492914 637954
rect 492294 637634 492914 637718
rect 492294 637398 492326 637634
rect 492562 637398 492646 637634
rect 492882 637398 492914 637634
rect 492294 601954 492914 637398
rect 492294 601718 492326 601954
rect 492562 601718 492646 601954
rect 492882 601718 492914 601954
rect 492294 601634 492914 601718
rect 492294 601398 492326 601634
rect 492562 601398 492646 601634
rect 492882 601398 492914 601634
rect 492294 565954 492914 601398
rect 492294 565718 492326 565954
rect 492562 565718 492646 565954
rect 492882 565718 492914 565954
rect 492294 565634 492914 565718
rect 492294 565398 492326 565634
rect 492562 565398 492646 565634
rect 492882 565398 492914 565634
rect 492294 529954 492914 565398
rect 492294 529718 492326 529954
rect 492562 529718 492646 529954
rect 492882 529718 492914 529954
rect 492294 529634 492914 529718
rect 492294 529398 492326 529634
rect 492562 529398 492646 529634
rect 492882 529398 492914 529634
rect 492294 493954 492914 529398
rect 492294 493718 492326 493954
rect 492562 493718 492646 493954
rect 492882 493718 492914 493954
rect 492294 493634 492914 493718
rect 492294 493398 492326 493634
rect 492562 493398 492646 493634
rect 492882 493398 492914 493634
rect 492294 457954 492914 493398
rect 492294 457718 492326 457954
rect 492562 457718 492646 457954
rect 492882 457718 492914 457954
rect 492294 457634 492914 457718
rect 492294 457398 492326 457634
rect 492562 457398 492646 457634
rect 492882 457398 492914 457634
rect 492294 421954 492914 457398
rect 492294 421718 492326 421954
rect 492562 421718 492646 421954
rect 492882 421718 492914 421954
rect 492294 421634 492914 421718
rect 492294 421398 492326 421634
rect 492562 421398 492646 421634
rect 492882 421398 492914 421634
rect 492294 385954 492914 421398
rect 492294 385718 492326 385954
rect 492562 385718 492646 385954
rect 492882 385718 492914 385954
rect 492294 385634 492914 385718
rect 492294 385398 492326 385634
rect 492562 385398 492646 385634
rect 492882 385398 492914 385634
rect 492294 349954 492914 385398
rect 492294 349718 492326 349954
rect 492562 349718 492646 349954
rect 492882 349718 492914 349954
rect 492294 349634 492914 349718
rect 492294 349398 492326 349634
rect 492562 349398 492646 349634
rect 492882 349398 492914 349634
rect 492294 313954 492914 349398
rect 492294 313718 492326 313954
rect 492562 313718 492646 313954
rect 492882 313718 492914 313954
rect 492294 313634 492914 313718
rect 492294 313398 492326 313634
rect 492562 313398 492646 313634
rect 492882 313398 492914 313634
rect 492294 277954 492914 313398
rect 492294 277718 492326 277954
rect 492562 277718 492646 277954
rect 492882 277718 492914 277954
rect 492294 277634 492914 277718
rect 492294 277398 492326 277634
rect 492562 277398 492646 277634
rect 492882 277398 492914 277634
rect 492294 241954 492914 277398
rect 492294 241718 492326 241954
rect 492562 241718 492646 241954
rect 492882 241718 492914 241954
rect 492294 241634 492914 241718
rect 492294 241398 492326 241634
rect 492562 241398 492646 241634
rect 492882 241398 492914 241634
rect 492294 205954 492914 241398
rect 492294 205718 492326 205954
rect 492562 205718 492646 205954
rect 492882 205718 492914 205954
rect 492294 205634 492914 205718
rect 492294 205398 492326 205634
rect 492562 205398 492646 205634
rect 492882 205398 492914 205634
rect 492294 169954 492914 205398
rect 492294 169718 492326 169954
rect 492562 169718 492646 169954
rect 492882 169718 492914 169954
rect 492294 169634 492914 169718
rect 492294 169398 492326 169634
rect 492562 169398 492646 169634
rect 492882 169398 492914 169634
rect 492294 133954 492914 169398
rect 492294 133718 492326 133954
rect 492562 133718 492646 133954
rect 492882 133718 492914 133954
rect 492294 133634 492914 133718
rect 492294 133398 492326 133634
rect 492562 133398 492646 133634
rect 492882 133398 492914 133634
rect 492294 97954 492914 133398
rect 492294 97718 492326 97954
rect 492562 97718 492646 97954
rect 492882 97718 492914 97954
rect 492294 97634 492914 97718
rect 492294 97398 492326 97634
rect 492562 97398 492646 97634
rect 492882 97398 492914 97634
rect 492294 61954 492914 97398
rect 492294 61718 492326 61954
rect 492562 61718 492646 61954
rect 492882 61718 492914 61954
rect 492294 61634 492914 61718
rect 492294 61398 492326 61634
rect 492562 61398 492646 61634
rect 492882 61398 492914 61634
rect 492294 25954 492914 61398
rect 492294 25718 492326 25954
rect 492562 25718 492646 25954
rect 492882 25718 492914 25954
rect 492294 25634 492914 25718
rect 492294 25398 492326 25634
rect 492562 25398 492646 25634
rect 492882 25398 492914 25634
rect 492294 -5146 492914 25398
rect 492294 -5382 492326 -5146
rect 492562 -5382 492646 -5146
rect 492882 -5382 492914 -5146
rect 492294 -5466 492914 -5382
rect 492294 -5702 492326 -5466
rect 492562 -5702 492646 -5466
rect 492882 -5702 492914 -5466
rect 492294 -7654 492914 -5702
rect 496794 710598 497414 711590
rect 496794 710362 496826 710598
rect 497062 710362 497146 710598
rect 497382 710362 497414 710598
rect 496794 710278 497414 710362
rect 496794 710042 496826 710278
rect 497062 710042 497146 710278
rect 497382 710042 497414 710278
rect 496794 678454 497414 710042
rect 496794 678218 496826 678454
rect 497062 678218 497146 678454
rect 497382 678218 497414 678454
rect 496794 678134 497414 678218
rect 496794 677898 496826 678134
rect 497062 677898 497146 678134
rect 497382 677898 497414 678134
rect 496794 642454 497414 677898
rect 496794 642218 496826 642454
rect 497062 642218 497146 642454
rect 497382 642218 497414 642454
rect 496794 642134 497414 642218
rect 496794 641898 496826 642134
rect 497062 641898 497146 642134
rect 497382 641898 497414 642134
rect 496794 606454 497414 641898
rect 496794 606218 496826 606454
rect 497062 606218 497146 606454
rect 497382 606218 497414 606454
rect 496794 606134 497414 606218
rect 496794 605898 496826 606134
rect 497062 605898 497146 606134
rect 497382 605898 497414 606134
rect 496794 570454 497414 605898
rect 496794 570218 496826 570454
rect 497062 570218 497146 570454
rect 497382 570218 497414 570454
rect 496794 570134 497414 570218
rect 496794 569898 496826 570134
rect 497062 569898 497146 570134
rect 497382 569898 497414 570134
rect 496794 534454 497414 569898
rect 496794 534218 496826 534454
rect 497062 534218 497146 534454
rect 497382 534218 497414 534454
rect 496794 534134 497414 534218
rect 496794 533898 496826 534134
rect 497062 533898 497146 534134
rect 497382 533898 497414 534134
rect 496794 498454 497414 533898
rect 496794 498218 496826 498454
rect 497062 498218 497146 498454
rect 497382 498218 497414 498454
rect 496794 498134 497414 498218
rect 496794 497898 496826 498134
rect 497062 497898 497146 498134
rect 497382 497898 497414 498134
rect 496794 462454 497414 497898
rect 496794 462218 496826 462454
rect 497062 462218 497146 462454
rect 497382 462218 497414 462454
rect 496794 462134 497414 462218
rect 496794 461898 496826 462134
rect 497062 461898 497146 462134
rect 497382 461898 497414 462134
rect 496794 426454 497414 461898
rect 496794 426218 496826 426454
rect 497062 426218 497146 426454
rect 497382 426218 497414 426454
rect 496794 426134 497414 426218
rect 496794 425898 496826 426134
rect 497062 425898 497146 426134
rect 497382 425898 497414 426134
rect 496794 390454 497414 425898
rect 496794 390218 496826 390454
rect 497062 390218 497146 390454
rect 497382 390218 497414 390454
rect 496794 390134 497414 390218
rect 496794 389898 496826 390134
rect 497062 389898 497146 390134
rect 497382 389898 497414 390134
rect 496794 354454 497414 389898
rect 496794 354218 496826 354454
rect 497062 354218 497146 354454
rect 497382 354218 497414 354454
rect 496794 354134 497414 354218
rect 496794 353898 496826 354134
rect 497062 353898 497146 354134
rect 497382 353898 497414 354134
rect 496794 318454 497414 353898
rect 496794 318218 496826 318454
rect 497062 318218 497146 318454
rect 497382 318218 497414 318454
rect 496794 318134 497414 318218
rect 496794 317898 496826 318134
rect 497062 317898 497146 318134
rect 497382 317898 497414 318134
rect 496794 282454 497414 317898
rect 496794 282218 496826 282454
rect 497062 282218 497146 282454
rect 497382 282218 497414 282454
rect 496794 282134 497414 282218
rect 496794 281898 496826 282134
rect 497062 281898 497146 282134
rect 497382 281898 497414 282134
rect 496794 246454 497414 281898
rect 496794 246218 496826 246454
rect 497062 246218 497146 246454
rect 497382 246218 497414 246454
rect 496794 246134 497414 246218
rect 496794 245898 496826 246134
rect 497062 245898 497146 246134
rect 497382 245898 497414 246134
rect 496794 210454 497414 245898
rect 496794 210218 496826 210454
rect 497062 210218 497146 210454
rect 497382 210218 497414 210454
rect 496794 210134 497414 210218
rect 496794 209898 496826 210134
rect 497062 209898 497146 210134
rect 497382 209898 497414 210134
rect 496794 174454 497414 209898
rect 496794 174218 496826 174454
rect 497062 174218 497146 174454
rect 497382 174218 497414 174454
rect 496794 174134 497414 174218
rect 496794 173898 496826 174134
rect 497062 173898 497146 174134
rect 497382 173898 497414 174134
rect 496794 138454 497414 173898
rect 496794 138218 496826 138454
rect 497062 138218 497146 138454
rect 497382 138218 497414 138454
rect 496794 138134 497414 138218
rect 496794 137898 496826 138134
rect 497062 137898 497146 138134
rect 497382 137898 497414 138134
rect 496794 102454 497414 137898
rect 496794 102218 496826 102454
rect 497062 102218 497146 102454
rect 497382 102218 497414 102454
rect 496794 102134 497414 102218
rect 496794 101898 496826 102134
rect 497062 101898 497146 102134
rect 497382 101898 497414 102134
rect 496794 66454 497414 101898
rect 496794 66218 496826 66454
rect 497062 66218 497146 66454
rect 497382 66218 497414 66454
rect 496794 66134 497414 66218
rect 496794 65898 496826 66134
rect 497062 65898 497146 66134
rect 497382 65898 497414 66134
rect 496794 30454 497414 65898
rect 496794 30218 496826 30454
rect 497062 30218 497146 30454
rect 497382 30218 497414 30454
rect 496794 30134 497414 30218
rect 496794 29898 496826 30134
rect 497062 29898 497146 30134
rect 497382 29898 497414 30134
rect 496794 -6106 497414 29898
rect 496794 -6342 496826 -6106
rect 497062 -6342 497146 -6106
rect 497382 -6342 497414 -6106
rect 496794 -6426 497414 -6342
rect 496794 -6662 496826 -6426
rect 497062 -6662 497146 -6426
rect 497382 -6662 497414 -6426
rect 496794 -7654 497414 -6662
rect 501294 711558 501914 711590
rect 501294 711322 501326 711558
rect 501562 711322 501646 711558
rect 501882 711322 501914 711558
rect 501294 711238 501914 711322
rect 501294 711002 501326 711238
rect 501562 711002 501646 711238
rect 501882 711002 501914 711238
rect 501294 682954 501914 711002
rect 501294 682718 501326 682954
rect 501562 682718 501646 682954
rect 501882 682718 501914 682954
rect 501294 682634 501914 682718
rect 501294 682398 501326 682634
rect 501562 682398 501646 682634
rect 501882 682398 501914 682634
rect 501294 646954 501914 682398
rect 501294 646718 501326 646954
rect 501562 646718 501646 646954
rect 501882 646718 501914 646954
rect 501294 646634 501914 646718
rect 501294 646398 501326 646634
rect 501562 646398 501646 646634
rect 501882 646398 501914 646634
rect 501294 610954 501914 646398
rect 501294 610718 501326 610954
rect 501562 610718 501646 610954
rect 501882 610718 501914 610954
rect 501294 610634 501914 610718
rect 501294 610398 501326 610634
rect 501562 610398 501646 610634
rect 501882 610398 501914 610634
rect 501294 574954 501914 610398
rect 501294 574718 501326 574954
rect 501562 574718 501646 574954
rect 501882 574718 501914 574954
rect 501294 574634 501914 574718
rect 501294 574398 501326 574634
rect 501562 574398 501646 574634
rect 501882 574398 501914 574634
rect 501294 538954 501914 574398
rect 501294 538718 501326 538954
rect 501562 538718 501646 538954
rect 501882 538718 501914 538954
rect 501294 538634 501914 538718
rect 501294 538398 501326 538634
rect 501562 538398 501646 538634
rect 501882 538398 501914 538634
rect 501294 502954 501914 538398
rect 501294 502718 501326 502954
rect 501562 502718 501646 502954
rect 501882 502718 501914 502954
rect 501294 502634 501914 502718
rect 501294 502398 501326 502634
rect 501562 502398 501646 502634
rect 501882 502398 501914 502634
rect 501294 466954 501914 502398
rect 501294 466718 501326 466954
rect 501562 466718 501646 466954
rect 501882 466718 501914 466954
rect 501294 466634 501914 466718
rect 501294 466398 501326 466634
rect 501562 466398 501646 466634
rect 501882 466398 501914 466634
rect 501294 430954 501914 466398
rect 501294 430718 501326 430954
rect 501562 430718 501646 430954
rect 501882 430718 501914 430954
rect 501294 430634 501914 430718
rect 501294 430398 501326 430634
rect 501562 430398 501646 430634
rect 501882 430398 501914 430634
rect 501294 394954 501914 430398
rect 501294 394718 501326 394954
rect 501562 394718 501646 394954
rect 501882 394718 501914 394954
rect 501294 394634 501914 394718
rect 501294 394398 501326 394634
rect 501562 394398 501646 394634
rect 501882 394398 501914 394634
rect 501294 358954 501914 394398
rect 501294 358718 501326 358954
rect 501562 358718 501646 358954
rect 501882 358718 501914 358954
rect 501294 358634 501914 358718
rect 501294 358398 501326 358634
rect 501562 358398 501646 358634
rect 501882 358398 501914 358634
rect 501294 322954 501914 358398
rect 501294 322718 501326 322954
rect 501562 322718 501646 322954
rect 501882 322718 501914 322954
rect 501294 322634 501914 322718
rect 501294 322398 501326 322634
rect 501562 322398 501646 322634
rect 501882 322398 501914 322634
rect 501294 286954 501914 322398
rect 501294 286718 501326 286954
rect 501562 286718 501646 286954
rect 501882 286718 501914 286954
rect 501294 286634 501914 286718
rect 501294 286398 501326 286634
rect 501562 286398 501646 286634
rect 501882 286398 501914 286634
rect 501294 250954 501914 286398
rect 501294 250718 501326 250954
rect 501562 250718 501646 250954
rect 501882 250718 501914 250954
rect 501294 250634 501914 250718
rect 501294 250398 501326 250634
rect 501562 250398 501646 250634
rect 501882 250398 501914 250634
rect 501294 214954 501914 250398
rect 501294 214718 501326 214954
rect 501562 214718 501646 214954
rect 501882 214718 501914 214954
rect 501294 214634 501914 214718
rect 501294 214398 501326 214634
rect 501562 214398 501646 214634
rect 501882 214398 501914 214634
rect 501294 178954 501914 214398
rect 501294 178718 501326 178954
rect 501562 178718 501646 178954
rect 501882 178718 501914 178954
rect 501294 178634 501914 178718
rect 501294 178398 501326 178634
rect 501562 178398 501646 178634
rect 501882 178398 501914 178634
rect 501294 142954 501914 178398
rect 501294 142718 501326 142954
rect 501562 142718 501646 142954
rect 501882 142718 501914 142954
rect 501294 142634 501914 142718
rect 501294 142398 501326 142634
rect 501562 142398 501646 142634
rect 501882 142398 501914 142634
rect 501294 106954 501914 142398
rect 501294 106718 501326 106954
rect 501562 106718 501646 106954
rect 501882 106718 501914 106954
rect 501294 106634 501914 106718
rect 501294 106398 501326 106634
rect 501562 106398 501646 106634
rect 501882 106398 501914 106634
rect 501294 70954 501914 106398
rect 501294 70718 501326 70954
rect 501562 70718 501646 70954
rect 501882 70718 501914 70954
rect 501294 70634 501914 70718
rect 501294 70398 501326 70634
rect 501562 70398 501646 70634
rect 501882 70398 501914 70634
rect 501294 34954 501914 70398
rect 501294 34718 501326 34954
rect 501562 34718 501646 34954
rect 501882 34718 501914 34954
rect 501294 34634 501914 34718
rect 501294 34398 501326 34634
rect 501562 34398 501646 34634
rect 501882 34398 501914 34634
rect 501294 -7066 501914 34398
rect 501294 -7302 501326 -7066
rect 501562 -7302 501646 -7066
rect 501882 -7302 501914 -7066
rect 501294 -7386 501914 -7302
rect 501294 -7622 501326 -7386
rect 501562 -7622 501646 -7386
rect 501882 -7622 501914 -7386
rect 501294 -7654 501914 -7622
rect 505794 704838 506414 711590
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 687454 506414 704282
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 505794 651454 506414 686898
rect 505794 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 506414 651454
rect 505794 651134 506414 651218
rect 505794 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 506414 651134
rect 505794 615454 506414 650898
rect 505794 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 506414 615454
rect 505794 615134 506414 615218
rect 505794 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 506414 615134
rect 505794 579454 506414 614898
rect 505794 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 506414 579454
rect 505794 579134 506414 579218
rect 505794 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 506414 579134
rect 505794 543454 506414 578898
rect 505794 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 506414 543454
rect 505794 543134 506414 543218
rect 505794 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 506414 543134
rect 505794 507454 506414 542898
rect 505794 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 506414 507454
rect 505794 507134 506414 507218
rect 505794 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 506414 507134
rect 505794 471454 506414 506898
rect 505794 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 506414 471454
rect 505794 471134 506414 471218
rect 505794 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 506414 471134
rect 505794 435454 506414 470898
rect 505794 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 506414 435454
rect 505794 435134 506414 435218
rect 505794 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 506414 435134
rect 505794 399454 506414 434898
rect 505794 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 506414 399454
rect 505794 399134 506414 399218
rect 505794 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 506414 399134
rect 505794 363454 506414 398898
rect 505794 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 506414 363454
rect 505794 363134 506414 363218
rect 505794 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 506414 363134
rect 505794 327454 506414 362898
rect 505794 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 506414 327454
rect 505794 327134 506414 327218
rect 505794 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 506414 327134
rect 505794 291454 506414 326898
rect 505794 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 506414 291454
rect 505794 291134 506414 291218
rect 505794 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 506414 291134
rect 505794 255454 506414 290898
rect 505794 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 506414 255454
rect 505794 255134 506414 255218
rect 505794 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 506414 255134
rect 505794 219454 506414 254898
rect 505794 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 506414 219454
rect 505794 219134 506414 219218
rect 505794 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 506414 219134
rect 505794 183454 506414 218898
rect 505794 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 506414 183454
rect 505794 183134 506414 183218
rect 505794 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 506414 183134
rect 505794 147454 506414 182898
rect 505794 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 506414 147454
rect 505794 147134 506414 147218
rect 505794 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 506414 147134
rect 505794 111454 506414 146898
rect 505794 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 506414 111454
rect 505794 111134 506414 111218
rect 505794 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 506414 111134
rect 505794 75454 506414 110898
rect 505794 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 506414 75454
rect 505794 75134 506414 75218
rect 505794 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 506414 75134
rect 505794 39454 506414 74898
rect 505794 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 506414 39454
rect 505794 39134 506414 39218
rect 505794 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 506414 39134
rect 505794 3454 506414 38898
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -7654 506414 -902
rect 510294 705798 510914 711590
rect 510294 705562 510326 705798
rect 510562 705562 510646 705798
rect 510882 705562 510914 705798
rect 510294 705478 510914 705562
rect 510294 705242 510326 705478
rect 510562 705242 510646 705478
rect 510882 705242 510914 705478
rect 510294 691954 510914 705242
rect 510294 691718 510326 691954
rect 510562 691718 510646 691954
rect 510882 691718 510914 691954
rect 510294 691634 510914 691718
rect 510294 691398 510326 691634
rect 510562 691398 510646 691634
rect 510882 691398 510914 691634
rect 510294 655954 510914 691398
rect 510294 655718 510326 655954
rect 510562 655718 510646 655954
rect 510882 655718 510914 655954
rect 510294 655634 510914 655718
rect 510294 655398 510326 655634
rect 510562 655398 510646 655634
rect 510882 655398 510914 655634
rect 510294 619954 510914 655398
rect 510294 619718 510326 619954
rect 510562 619718 510646 619954
rect 510882 619718 510914 619954
rect 510294 619634 510914 619718
rect 510294 619398 510326 619634
rect 510562 619398 510646 619634
rect 510882 619398 510914 619634
rect 510294 583954 510914 619398
rect 510294 583718 510326 583954
rect 510562 583718 510646 583954
rect 510882 583718 510914 583954
rect 510294 583634 510914 583718
rect 510294 583398 510326 583634
rect 510562 583398 510646 583634
rect 510882 583398 510914 583634
rect 510294 547954 510914 583398
rect 510294 547718 510326 547954
rect 510562 547718 510646 547954
rect 510882 547718 510914 547954
rect 510294 547634 510914 547718
rect 510294 547398 510326 547634
rect 510562 547398 510646 547634
rect 510882 547398 510914 547634
rect 510294 511954 510914 547398
rect 510294 511718 510326 511954
rect 510562 511718 510646 511954
rect 510882 511718 510914 511954
rect 510294 511634 510914 511718
rect 510294 511398 510326 511634
rect 510562 511398 510646 511634
rect 510882 511398 510914 511634
rect 510294 475954 510914 511398
rect 510294 475718 510326 475954
rect 510562 475718 510646 475954
rect 510882 475718 510914 475954
rect 510294 475634 510914 475718
rect 510294 475398 510326 475634
rect 510562 475398 510646 475634
rect 510882 475398 510914 475634
rect 510294 439954 510914 475398
rect 510294 439718 510326 439954
rect 510562 439718 510646 439954
rect 510882 439718 510914 439954
rect 510294 439634 510914 439718
rect 510294 439398 510326 439634
rect 510562 439398 510646 439634
rect 510882 439398 510914 439634
rect 510294 403954 510914 439398
rect 510294 403718 510326 403954
rect 510562 403718 510646 403954
rect 510882 403718 510914 403954
rect 510294 403634 510914 403718
rect 510294 403398 510326 403634
rect 510562 403398 510646 403634
rect 510882 403398 510914 403634
rect 510294 367954 510914 403398
rect 510294 367718 510326 367954
rect 510562 367718 510646 367954
rect 510882 367718 510914 367954
rect 510294 367634 510914 367718
rect 510294 367398 510326 367634
rect 510562 367398 510646 367634
rect 510882 367398 510914 367634
rect 510294 331954 510914 367398
rect 510294 331718 510326 331954
rect 510562 331718 510646 331954
rect 510882 331718 510914 331954
rect 510294 331634 510914 331718
rect 510294 331398 510326 331634
rect 510562 331398 510646 331634
rect 510882 331398 510914 331634
rect 510294 295954 510914 331398
rect 510294 295718 510326 295954
rect 510562 295718 510646 295954
rect 510882 295718 510914 295954
rect 510294 295634 510914 295718
rect 510294 295398 510326 295634
rect 510562 295398 510646 295634
rect 510882 295398 510914 295634
rect 510294 259954 510914 295398
rect 510294 259718 510326 259954
rect 510562 259718 510646 259954
rect 510882 259718 510914 259954
rect 510294 259634 510914 259718
rect 510294 259398 510326 259634
rect 510562 259398 510646 259634
rect 510882 259398 510914 259634
rect 510294 223954 510914 259398
rect 510294 223718 510326 223954
rect 510562 223718 510646 223954
rect 510882 223718 510914 223954
rect 510294 223634 510914 223718
rect 510294 223398 510326 223634
rect 510562 223398 510646 223634
rect 510882 223398 510914 223634
rect 510294 187954 510914 223398
rect 510294 187718 510326 187954
rect 510562 187718 510646 187954
rect 510882 187718 510914 187954
rect 510294 187634 510914 187718
rect 510294 187398 510326 187634
rect 510562 187398 510646 187634
rect 510882 187398 510914 187634
rect 510294 151954 510914 187398
rect 510294 151718 510326 151954
rect 510562 151718 510646 151954
rect 510882 151718 510914 151954
rect 510294 151634 510914 151718
rect 510294 151398 510326 151634
rect 510562 151398 510646 151634
rect 510882 151398 510914 151634
rect 510294 115954 510914 151398
rect 510294 115718 510326 115954
rect 510562 115718 510646 115954
rect 510882 115718 510914 115954
rect 510294 115634 510914 115718
rect 510294 115398 510326 115634
rect 510562 115398 510646 115634
rect 510882 115398 510914 115634
rect 510294 79954 510914 115398
rect 510294 79718 510326 79954
rect 510562 79718 510646 79954
rect 510882 79718 510914 79954
rect 510294 79634 510914 79718
rect 510294 79398 510326 79634
rect 510562 79398 510646 79634
rect 510882 79398 510914 79634
rect 510294 43954 510914 79398
rect 510294 43718 510326 43954
rect 510562 43718 510646 43954
rect 510882 43718 510914 43954
rect 510294 43634 510914 43718
rect 510294 43398 510326 43634
rect 510562 43398 510646 43634
rect 510882 43398 510914 43634
rect 510294 7954 510914 43398
rect 510294 7718 510326 7954
rect 510562 7718 510646 7954
rect 510882 7718 510914 7954
rect 510294 7634 510914 7718
rect 510294 7398 510326 7634
rect 510562 7398 510646 7634
rect 510882 7398 510914 7634
rect 510294 -1306 510914 7398
rect 510294 -1542 510326 -1306
rect 510562 -1542 510646 -1306
rect 510882 -1542 510914 -1306
rect 510294 -1626 510914 -1542
rect 510294 -1862 510326 -1626
rect 510562 -1862 510646 -1626
rect 510882 -1862 510914 -1626
rect 510294 -7654 510914 -1862
rect 514794 706758 515414 711590
rect 514794 706522 514826 706758
rect 515062 706522 515146 706758
rect 515382 706522 515414 706758
rect 514794 706438 515414 706522
rect 514794 706202 514826 706438
rect 515062 706202 515146 706438
rect 515382 706202 515414 706438
rect 514794 696454 515414 706202
rect 514794 696218 514826 696454
rect 515062 696218 515146 696454
rect 515382 696218 515414 696454
rect 514794 696134 515414 696218
rect 514794 695898 514826 696134
rect 515062 695898 515146 696134
rect 515382 695898 515414 696134
rect 514794 660454 515414 695898
rect 514794 660218 514826 660454
rect 515062 660218 515146 660454
rect 515382 660218 515414 660454
rect 514794 660134 515414 660218
rect 514794 659898 514826 660134
rect 515062 659898 515146 660134
rect 515382 659898 515414 660134
rect 514794 624454 515414 659898
rect 514794 624218 514826 624454
rect 515062 624218 515146 624454
rect 515382 624218 515414 624454
rect 514794 624134 515414 624218
rect 514794 623898 514826 624134
rect 515062 623898 515146 624134
rect 515382 623898 515414 624134
rect 514794 588454 515414 623898
rect 514794 588218 514826 588454
rect 515062 588218 515146 588454
rect 515382 588218 515414 588454
rect 514794 588134 515414 588218
rect 514794 587898 514826 588134
rect 515062 587898 515146 588134
rect 515382 587898 515414 588134
rect 514794 552454 515414 587898
rect 514794 552218 514826 552454
rect 515062 552218 515146 552454
rect 515382 552218 515414 552454
rect 514794 552134 515414 552218
rect 514794 551898 514826 552134
rect 515062 551898 515146 552134
rect 515382 551898 515414 552134
rect 514794 516454 515414 551898
rect 514794 516218 514826 516454
rect 515062 516218 515146 516454
rect 515382 516218 515414 516454
rect 514794 516134 515414 516218
rect 514794 515898 514826 516134
rect 515062 515898 515146 516134
rect 515382 515898 515414 516134
rect 514794 480454 515414 515898
rect 514794 480218 514826 480454
rect 515062 480218 515146 480454
rect 515382 480218 515414 480454
rect 514794 480134 515414 480218
rect 514794 479898 514826 480134
rect 515062 479898 515146 480134
rect 515382 479898 515414 480134
rect 514794 444454 515414 479898
rect 514794 444218 514826 444454
rect 515062 444218 515146 444454
rect 515382 444218 515414 444454
rect 514794 444134 515414 444218
rect 514794 443898 514826 444134
rect 515062 443898 515146 444134
rect 515382 443898 515414 444134
rect 514794 408454 515414 443898
rect 514794 408218 514826 408454
rect 515062 408218 515146 408454
rect 515382 408218 515414 408454
rect 514794 408134 515414 408218
rect 514794 407898 514826 408134
rect 515062 407898 515146 408134
rect 515382 407898 515414 408134
rect 514794 372454 515414 407898
rect 514794 372218 514826 372454
rect 515062 372218 515146 372454
rect 515382 372218 515414 372454
rect 514794 372134 515414 372218
rect 514794 371898 514826 372134
rect 515062 371898 515146 372134
rect 515382 371898 515414 372134
rect 514794 336454 515414 371898
rect 514794 336218 514826 336454
rect 515062 336218 515146 336454
rect 515382 336218 515414 336454
rect 514794 336134 515414 336218
rect 514794 335898 514826 336134
rect 515062 335898 515146 336134
rect 515382 335898 515414 336134
rect 514794 300454 515414 335898
rect 514794 300218 514826 300454
rect 515062 300218 515146 300454
rect 515382 300218 515414 300454
rect 514794 300134 515414 300218
rect 514794 299898 514826 300134
rect 515062 299898 515146 300134
rect 515382 299898 515414 300134
rect 514794 264454 515414 299898
rect 514794 264218 514826 264454
rect 515062 264218 515146 264454
rect 515382 264218 515414 264454
rect 514794 264134 515414 264218
rect 514794 263898 514826 264134
rect 515062 263898 515146 264134
rect 515382 263898 515414 264134
rect 514794 228454 515414 263898
rect 514794 228218 514826 228454
rect 515062 228218 515146 228454
rect 515382 228218 515414 228454
rect 514794 228134 515414 228218
rect 514794 227898 514826 228134
rect 515062 227898 515146 228134
rect 515382 227898 515414 228134
rect 514794 192454 515414 227898
rect 514794 192218 514826 192454
rect 515062 192218 515146 192454
rect 515382 192218 515414 192454
rect 514794 192134 515414 192218
rect 514794 191898 514826 192134
rect 515062 191898 515146 192134
rect 515382 191898 515414 192134
rect 514794 156454 515414 191898
rect 514794 156218 514826 156454
rect 515062 156218 515146 156454
rect 515382 156218 515414 156454
rect 514794 156134 515414 156218
rect 514794 155898 514826 156134
rect 515062 155898 515146 156134
rect 515382 155898 515414 156134
rect 514794 120454 515414 155898
rect 514794 120218 514826 120454
rect 515062 120218 515146 120454
rect 515382 120218 515414 120454
rect 514794 120134 515414 120218
rect 514794 119898 514826 120134
rect 515062 119898 515146 120134
rect 515382 119898 515414 120134
rect 514794 84454 515414 119898
rect 514794 84218 514826 84454
rect 515062 84218 515146 84454
rect 515382 84218 515414 84454
rect 514794 84134 515414 84218
rect 514794 83898 514826 84134
rect 515062 83898 515146 84134
rect 515382 83898 515414 84134
rect 514794 48454 515414 83898
rect 514794 48218 514826 48454
rect 515062 48218 515146 48454
rect 515382 48218 515414 48454
rect 514794 48134 515414 48218
rect 514794 47898 514826 48134
rect 515062 47898 515146 48134
rect 515382 47898 515414 48134
rect 514794 12454 515414 47898
rect 514794 12218 514826 12454
rect 515062 12218 515146 12454
rect 515382 12218 515414 12454
rect 514794 12134 515414 12218
rect 514794 11898 514826 12134
rect 515062 11898 515146 12134
rect 515382 11898 515414 12134
rect 514794 -2266 515414 11898
rect 514794 -2502 514826 -2266
rect 515062 -2502 515146 -2266
rect 515382 -2502 515414 -2266
rect 514794 -2586 515414 -2502
rect 514794 -2822 514826 -2586
rect 515062 -2822 515146 -2586
rect 515382 -2822 515414 -2586
rect 514794 -7654 515414 -2822
rect 519294 707718 519914 711590
rect 519294 707482 519326 707718
rect 519562 707482 519646 707718
rect 519882 707482 519914 707718
rect 519294 707398 519914 707482
rect 519294 707162 519326 707398
rect 519562 707162 519646 707398
rect 519882 707162 519914 707398
rect 519294 700954 519914 707162
rect 519294 700718 519326 700954
rect 519562 700718 519646 700954
rect 519882 700718 519914 700954
rect 519294 700634 519914 700718
rect 519294 700398 519326 700634
rect 519562 700398 519646 700634
rect 519882 700398 519914 700634
rect 519294 664954 519914 700398
rect 519294 664718 519326 664954
rect 519562 664718 519646 664954
rect 519882 664718 519914 664954
rect 519294 664634 519914 664718
rect 519294 664398 519326 664634
rect 519562 664398 519646 664634
rect 519882 664398 519914 664634
rect 519294 628954 519914 664398
rect 519294 628718 519326 628954
rect 519562 628718 519646 628954
rect 519882 628718 519914 628954
rect 519294 628634 519914 628718
rect 519294 628398 519326 628634
rect 519562 628398 519646 628634
rect 519882 628398 519914 628634
rect 519294 592954 519914 628398
rect 519294 592718 519326 592954
rect 519562 592718 519646 592954
rect 519882 592718 519914 592954
rect 519294 592634 519914 592718
rect 519294 592398 519326 592634
rect 519562 592398 519646 592634
rect 519882 592398 519914 592634
rect 519294 556954 519914 592398
rect 519294 556718 519326 556954
rect 519562 556718 519646 556954
rect 519882 556718 519914 556954
rect 519294 556634 519914 556718
rect 519294 556398 519326 556634
rect 519562 556398 519646 556634
rect 519882 556398 519914 556634
rect 519294 520954 519914 556398
rect 519294 520718 519326 520954
rect 519562 520718 519646 520954
rect 519882 520718 519914 520954
rect 519294 520634 519914 520718
rect 519294 520398 519326 520634
rect 519562 520398 519646 520634
rect 519882 520398 519914 520634
rect 519294 484954 519914 520398
rect 519294 484718 519326 484954
rect 519562 484718 519646 484954
rect 519882 484718 519914 484954
rect 519294 484634 519914 484718
rect 519294 484398 519326 484634
rect 519562 484398 519646 484634
rect 519882 484398 519914 484634
rect 519294 448954 519914 484398
rect 519294 448718 519326 448954
rect 519562 448718 519646 448954
rect 519882 448718 519914 448954
rect 519294 448634 519914 448718
rect 519294 448398 519326 448634
rect 519562 448398 519646 448634
rect 519882 448398 519914 448634
rect 519294 412954 519914 448398
rect 519294 412718 519326 412954
rect 519562 412718 519646 412954
rect 519882 412718 519914 412954
rect 519294 412634 519914 412718
rect 519294 412398 519326 412634
rect 519562 412398 519646 412634
rect 519882 412398 519914 412634
rect 519294 376954 519914 412398
rect 519294 376718 519326 376954
rect 519562 376718 519646 376954
rect 519882 376718 519914 376954
rect 519294 376634 519914 376718
rect 519294 376398 519326 376634
rect 519562 376398 519646 376634
rect 519882 376398 519914 376634
rect 519294 340954 519914 376398
rect 519294 340718 519326 340954
rect 519562 340718 519646 340954
rect 519882 340718 519914 340954
rect 519294 340634 519914 340718
rect 519294 340398 519326 340634
rect 519562 340398 519646 340634
rect 519882 340398 519914 340634
rect 519294 304954 519914 340398
rect 519294 304718 519326 304954
rect 519562 304718 519646 304954
rect 519882 304718 519914 304954
rect 519294 304634 519914 304718
rect 519294 304398 519326 304634
rect 519562 304398 519646 304634
rect 519882 304398 519914 304634
rect 519294 268954 519914 304398
rect 519294 268718 519326 268954
rect 519562 268718 519646 268954
rect 519882 268718 519914 268954
rect 519294 268634 519914 268718
rect 519294 268398 519326 268634
rect 519562 268398 519646 268634
rect 519882 268398 519914 268634
rect 519294 232954 519914 268398
rect 519294 232718 519326 232954
rect 519562 232718 519646 232954
rect 519882 232718 519914 232954
rect 519294 232634 519914 232718
rect 519294 232398 519326 232634
rect 519562 232398 519646 232634
rect 519882 232398 519914 232634
rect 519294 196954 519914 232398
rect 519294 196718 519326 196954
rect 519562 196718 519646 196954
rect 519882 196718 519914 196954
rect 519294 196634 519914 196718
rect 519294 196398 519326 196634
rect 519562 196398 519646 196634
rect 519882 196398 519914 196634
rect 519294 160954 519914 196398
rect 519294 160718 519326 160954
rect 519562 160718 519646 160954
rect 519882 160718 519914 160954
rect 519294 160634 519914 160718
rect 519294 160398 519326 160634
rect 519562 160398 519646 160634
rect 519882 160398 519914 160634
rect 519294 124954 519914 160398
rect 519294 124718 519326 124954
rect 519562 124718 519646 124954
rect 519882 124718 519914 124954
rect 519294 124634 519914 124718
rect 519294 124398 519326 124634
rect 519562 124398 519646 124634
rect 519882 124398 519914 124634
rect 519294 88954 519914 124398
rect 519294 88718 519326 88954
rect 519562 88718 519646 88954
rect 519882 88718 519914 88954
rect 519294 88634 519914 88718
rect 519294 88398 519326 88634
rect 519562 88398 519646 88634
rect 519882 88398 519914 88634
rect 519294 52954 519914 88398
rect 519294 52718 519326 52954
rect 519562 52718 519646 52954
rect 519882 52718 519914 52954
rect 519294 52634 519914 52718
rect 519294 52398 519326 52634
rect 519562 52398 519646 52634
rect 519882 52398 519914 52634
rect 519294 16954 519914 52398
rect 519294 16718 519326 16954
rect 519562 16718 519646 16954
rect 519882 16718 519914 16954
rect 519294 16634 519914 16718
rect 519294 16398 519326 16634
rect 519562 16398 519646 16634
rect 519882 16398 519914 16634
rect 519294 -3226 519914 16398
rect 519294 -3462 519326 -3226
rect 519562 -3462 519646 -3226
rect 519882 -3462 519914 -3226
rect 519294 -3546 519914 -3462
rect 519294 -3782 519326 -3546
rect 519562 -3782 519646 -3546
rect 519882 -3782 519914 -3546
rect 519294 -7654 519914 -3782
rect 523794 708678 524414 711590
rect 523794 708442 523826 708678
rect 524062 708442 524146 708678
rect 524382 708442 524414 708678
rect 523794 708358 524414 708442
rect 523794 708122 523826 708358
rect 524062 708122 524146 708358
rect 524382 708122 524414 708358
rect 523794 669454 524414 708122
rect 523794 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 524414 669454
rect 523794 669134 524414 669218
rect 523794 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 524414 669134
rect 523794 633454 524414 668898
rect 523794 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 524414 633454
rect 523794 633134 524414 633218
rect 523794 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 524414 633134
rect 523794 597454 524414 632898
rect 523794 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 524414 597454
rect 523794 597134 524414 597218
rect 523794 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 524414 597134
rect 523794 561454 524414 596898
rect 523794 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 524414 561454
rect 523794 561134 524414 561218
rect 523794 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 524414 561134
rect 523794 525454 524414 560898
rect 523794 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 524414 525454
rect 523794 525134 524414 525218
rect 523794 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 524414 525134
rect 523794 489454 524414 524898
rect 523794 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 524414 489454
rect 523794 489134 524414 489218
rect 523794 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 524414 489134
rect 523794 453454 524414 488898
rect 523794 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 524414 453454
rect 523794 453134 524414 453218
rect 523794 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 524414 453134
rect 523794 417454 524414 452898
rect 523794 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 524414 417454
rect 523794 417134 524414 417218
rect 523794 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 524414 417134
rect 523794 381454 524414 416898
rect 523794 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 524414 381454
rect 523794 381134 524414 381218
rect 523794 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 524414 381134
rect 523794 345454 524414 380898
rect 523794 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 524414 345454
rect 523794 345134 524414 345218
rect 523794 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 524414 345134
rect 523794 309454 524414 344898
rect 523794 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 524414 309454
rect 523794 309134 524414 309218
rect 523794 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 524414 309134
rect 523794 273454 524414 308898
rect 523794 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 524414 273454
rect 523794 273134 524414 273218
rect 523794 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 524414 273134
rect 523794 237454 524414 272898
rect 523794 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 524414 237454
rect 523794 237134 524414 237218
rect 523794 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 524414 237134
rect 523794 201454 524414 236898
rect 523794 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 524414 201454
rect 523794 201134 524414 201218
rect 523794 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 524414 201134
rect 523794 165454 524414 200898
rect 523794 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 524414 165454
rect 523794 165134 524414 165218
rect 523794 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 524414 165134
rect 523794 129454 524414 164898
rect 523794 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 524414 129454
rect 523794 129134 524414 129218
rect 523794 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 524414 129134
rect 523794 93454 524414 128898
rect 523794 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 524414 93454
rect 523794 93134 524414 93218
rect 523794 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 524414 93134
rect 523794 57454 524414 92898
rect 523794 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 524414 57454
rect 523794 57134 524414 57218
rect 523794 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 524414 57134
rect 523794 21454 524414 56898
rect 523794 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 524414 21454
rect 523794 21134 524414 21218
rect 523794 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 524414 21134
rect 523794 -4186 524414 20898
rect 523794 -4422 523826 -4186
rect 524062 -4422 524146 -4186
rect 524382 -4422 524414 -4186
rect 523794 -4506 524414 -4422
rect 523794 -4742 523826 -4506
rect 524062 -4742 524146 -4506
rect 524382 -4742 524414 -4506
rect 523794 -7654 524414 -4742
rect 528294 709638 528914 711590
rect 528294 709402 528326 709638
rect 528562 709402 528646 709638
rect 528882 709402 528914 709638
rect 528294 709318 528914 709402
rect 528294 709082 528326 709318
rect 528562 709082 528646 709318
rect 528882 709082 528914 709318
rect 528294 673954 528914 709082
rect 528294 673718 528326 673954
rect 528562 673718 528646 673954
rect 528882 673718 528914 673954
rect 528294 673634 528914 673718
rect 528294 673398 528326 673634
rect 528562 673398 528646 673634
rect 528882 673398 528914 673634
rect 528294 637954 528914 673398
rect 528294 637718 528326 637954
rect 528562 637718 528646 637954
rect 528882 637718 528914 637954
rect 528294 637634 528914 637718
rect 528294 637398 528326 637634
rect 528562 637398 528646 637634
rect 528882 637398 528914 637634
rect 528294 601954 528914 637398
rect 528294 601718 528326 601954
rect 528562 601718 528646 601954
rect 528882 601718 528914 601954
rect 528294 601634 528914 601718
rect 528294 601398 528326 601634
rect 528562 601398 528646 601634
rect 528882 601398 528914 601634
rect 528294 565954 528914 601398
rect 528294 565718 528326 565954
rect 528562 565718 528646 565954
rect 528882 565718 528914 565954
rect 528294 565634 528914 565718
rect 528294 565398 528326 565634
rect 528562 565398 528646 565634
rect 528882 565398 528914 565634
rect 528294 529954 528914 565398
rect 528294 529718 528326 529954
rect 528562 529718 528646 529954
rect 528882 529718 528914 529954
rect 528294 529634 528914 529718
rect 528294 529398 528326 529634
rect 528562 529398 528646 529634
rect 528882 529398 528914 529634
rect 528294 493954 528914 529398
rect 528294 493718 528326 493954
rect 528562 493718 528646 493954
rect 528882 493718 528914 493954
rect 528294 493634 528914 493718
rect 528294 493398 528326 493634
rect 528562 493398 528646 493634
rect 528882 493398 528914 493634
rect 528294 457954 528914 493398
rect 528294 457718 528326 457954
rect 528562 457718 528646 457954
rect 528882 457718 528914 457954
rect 528294 457634 528914 457718
rect 528294 457398 528326 457634
rect 528562 457398 528646 457634
rect 528882 457398 528914 457634
rect 528294 421954 528914 457398
rect 528294 421718 528326 421954
rect 528562 421718 528646 421954
rect 528882 421718 528914 421954
rect 528294 421634 528914 421718
rect 528294 421398 528326 421634
rect 528562 421398 528646 421634
rect 528882 421398 528914 421634
rect 528294 385954 528914 421398
rect 528294 385718 528326 385954
rect 528562 385718 528646 385954
rect 528882 385718 528914 385954
rect 528294 385634 528914 385718
rect 528294 385398 528326 385634
rect 528562 385398 528646 385634
rect 528882 385398 528914 385634
rect 528294 349954 528914 385398
rect 528294 349718 528326 349954
rect 528562 349718 528646 349954
rect 528882 349718 528914 349954
rect 528294 349634 528914 349718
rect 528294 349398 528326 349634
rect 528562 349398 528646 349634
rect 528882 349398 528914 349634
rect 528294 313954 528914 349398
rect 528294 313718 528326 313954
rect 528562 313718 528646 313954
rect 528882 313718 528914 313954
rect 528294 313634 528914 313718
rect 528294 313398 528326 313634
rect 528562 313398 528646 313634
rect 528882 313398 528914 313634
rect 528294 277954 528914 313398
rect 528294 277718 528326 277954
rect 528562 277718 528646 277954
rect 528882 277718 528914 277954
rect 528294 277634 528914 277718
rect 528294 277398 528326 277634
rect 528562 277398 528646 277634
rect 528882 277398 528914 277634
rect 528294 241954 528914 277398
rect 528294 241718 528326 241954
rect 528562 241718 528646 241954
rect 528882 241718 528914 241954
rect 528294 241634 528914 241718
rect 528294 241398 528326 241634
rect 528562 241398 528646 241634
rect 528882 241398 528914 241634
rect 528294 205954 528914 241398
rect 528294 205718 528326 205954
rect 528562 205718 528646 205954
rect 528882 205718 528914 205954
rect 528294 205634 528914 205718
rect 528294 205398 528326 205634
rect 528562 205398 528646 205634
rect 528882 205398 528914 205634
rect 528294 169954 528914 205398
rect 528294 169718 528326 169954
rect 528562 169718 528646 169954
rect 528882 169718 528914 169954
rect 528294 169634 528914 169718
rect 528294 169398 528326 169634
rect 528562 169398 528646 169634
rect 528882 169398 528914 169634
rect 528294 133954 528914 169398
rect 528294 133718 528326 133954
rect 528562 133718 528646 133954
rect 528882 133718 528914 133954
rect 528294 133634 528914 133718
rect 528294 133398 528326 133634
rect 528562 133398 528646 133634
rect 528882 133398 528914 133634
rect 528294 97954 528914 133398
rect 528294 97718 528326 97954
rect 528562 97718 528646 97954
rect 528882 97718 528914 97954
rect 528294 97634 528914 97718
rect 528294 97398 528326 97634
rect 528562 97398 528646 97634
rect 528882 97398 528914 97634
rect 528294 61954 528914 97398
rect 528294 61718 528326 61954
rect 528562 61718 528646 61954
rect 528882 61718 528914 61954
rect 528294 61634 528914 61718
rect 528294 61398 528326 61634
rect 528562 61398 528646 61634
rect 528882 61398 528914 61634
rect 528294 25954 528914 61398
rect 528294 25718 528326 25954
rect 528562 25718 528646 25954
rect 528882 25718 528914 25954
rect 528294 25634 528914 25718
rect 528294 25398 528326 25634
rect 528562 25398 528646 25634
rect 528882 25398 528914 25634
rect 528294 -5146 528914 25398
rect 528294 -5382 528326 -5146
rect 528562 -5382 528646 -5146
rect 528882 -5382 528914 -5146
rect 528294 -5466 528914 -5382
rect 528294 -5702 528326 -5466
rect 528562 -5702 528646 -5466
rect 528882 -5702 528914 -5466
rect 528294 -7654 528914 -5702
rect 532794 710598 533414 711590
rect 532794 710362 532826 710598
rect 533062 710362 533146 710598
rect 533382 710362 533414 710598
rect 532794 710278 533414 710362
rect 532794 710042 532826 710278
rect 533062 710042 533146 710278
rect 533382 710042 533414 710278
rect 532794 678454 533414 710042
rect 532794 678218 532826 678454
rect 533062 678218 533146 678454
rect 533382 678218 533414 678454
rect 532794 678134 533414 678218
rect 532794 677898 532826 678134
rect 533062 677898 533146 678134
rect 533382 677898 533414 678134
rect 532794 642454 533414 677898
rect 532794 642218 532826 642454
rect 533062 642218 533146 642454
rect 533382 642218 533414 642454
rect 532794 642134 533414 642218
rect 532794 641898 532826 642134
rect 533062 641898 533146 642134
rect 533382 641898 533414 642134
rect 532794 606454 533414 641898
rect 532794 606218 532826 606454
rect 533062 606218 533146 606454
rect 533382 606218 533414 606454
rect 532794 606134 533414 606218
rect 532794 605898 532826 606134
rect 533062 605898 533146 606134
rect 533382 605898 533414 606134
rect 532794 570454 533414 605898
rect 532794 570218 532826 570454
rect 533062 570218 533146 570454
rect 533382 570218 533414 570454
rect 532794 570134 533414 570218
rect 532794 569898 532826 570134
rect 533062 569898 533146 570134
rect 533382 569898 533414 570134
rect 532794 534454 533414 569898
rect 532794 534218 532826 534454
rect 533062 534218 533146 534454
rect 533382 534218 533414 534454
rect 532794 534134 533414 534218
rect 532794 533898 532826 534134
rect 533062 533898 533146 534134
rect 533382 533898 533414 534134
rect 532794 498454 533414 533898
rect 532794 498218 532826 498454
rect 533062 498218 533146 498454
rect 533382 498218 533414 498454
rect 532794 498134 533414 498218
rect 532794 497898 532826 498134
rect 533062 497898 533146 498134
rect 533382 497898 533414 498134
rect 532794 462454 533414 497898
rect 532794 462218 532826 462454
rect 533062 462218 533146 462454
rect 533382 462218 533414 462454
rect 532794 462134 533414 462218
rect 532794 461898 532826 462134
rect 533062 461898 533146 462134
rect 533382 461898 533414 462134
rect 532794 426454 533414 461898
rect 532794 426218 532826 426454
rect 533062 426218 533146 426454
rect 533382 426218 533414 426454
rect 532794 426134 533414 426218
rect 532794 425898 532826 426134
rect 533062 425898 533146 426134
rect 533382 425898 533414 426134
rect 532794 390454 533414 425898
rect 532794 390218 532826 390454
rect 533062 390218 533146 390454
rect 533382 390218 533414 390454
rect 532794 390134 533414 390218
rect 532794 389898 532826 390134
rect 533062 389898 533146 390134
rect 533382 389898 533414 390134
rect 532794 354454 533414 389898
rect 532794 354218 532826 354454
rect 533062 354218 533146 354454
rect 533382 354218 533414 354454
rect 532794 354134 533414 354218
rect 532794 353898 532826 354134
rect 533062 353898 533146 354134
rect 533382 353898 533414 354134
rect 532794 318454 533414 353898
rect 532794 318218 532826 318454
rect 533062 318218 533146 318454
rect 533382 318218 533414 318454
rect 532794 318134 533414 318218
rect 532794 317898 532826 318134
rect 533062 317898 533146 318134
rect 533382 317898 533414 318134
rect 532794 282454 533414 317898
rect 532794 282218 532826 282454
rect 533062 282218 533146 282454
rect 533382 282218 533414 282454
rect 532794 282134 533414 282218
rect 532794 281898 532826 282134
rect 533062 281898 533146 282134
rect 533382 281898 533414 282134
rect 532794 246454 533414 281898
rect 532794 246218 532826 246454
rect 533062 246218 533146 246454
rect 533382 246218 533414 246454
rect 532794 246134 533414 246218
rect 532794 245898 532826 246134
rect 533062 245898 533146 246134
rect 533382 245898 533414 246134
rect 532794 210454 533414 245898
rect 532794 210218 532826 210454
rect 533062 210218 533146 210454
rect 533382 210218 533414 210454
rect 532794 210134 533414 210218
rect 532794 209898 532826 210134
rect 533062 209898 533146 210134
rect 533382 209898 533414 210134
rect 532794 174454 533414 209898
rect 532794 174218 532826 174454
rect 533062 174218 533146 174454
rect 533382 174218 533414 174454
rect 532794 174134 533414 174218
rect 532794 173898 532826 174134
rect 533062 173898 533146 174134
rect 533382 173898 533414 174134
rect 532794 138454 533414 173898
rect 532794 138218 532826 138454
rect 533062 138218 533146 138454
rect 533382 138218 533414 138454
rect 532794 138134 533414 138218
rect 532794 137898 532826 138134
rect 533062 137898 533146 138134
rect 533382 137898 533414 138134
rect 532794 102454 533414 137898
rect 532794 102218 532826 102454
rect 533062 102218 533146 102454
rect 533382 102218 533414 102454
rect 532794 102134 533414 102218
rect 532794 101898 532826 102134
rect 533062 101898 533146 102134
rect 533382 101898 533414 102134
rect 532794 66454 533414 101898
rect 532794 66218 532826 66454
rect 533062 66218 533146 66454
rect 533382 66218 533414 66454
rect 532794 66134 533414 66218
rect 532794 65898 532826 66134
rect 533062 65898 533146 66134
rect 533382 65898 533414 66134
rect 532794 30454 533414 65898
rect 532794 30218 532826 30454
rect 533062 30218 533146 30454
rect 533382 30218 533414 30454
rect 532794 30134 533414 30218
rect 532794 29898 532826 30134
rect 533062 29898 533146 30134
rect 533382 29898 533414 30134
rect 532794 -6106 533414 29898
rect 532794 -6342 532826 -6106
rect 533062 -6342 533146 -6106
rect 533382 -6342 533414 -6106
rect 532794 -6426 533414 -6342
rect 532794 -6662 532826 -6426
rect 533062 -6662 533146 -6426
rect 533382 -6662 533414 -6426
rect 532794 -7654 533414 -6662
rect 537294 711558 537914 711590
rect 537294 711322 537326 711558
rect 537562 711322 537646 711558
rect 537882 711322 537914 711558
rect 537294 711238 537914 711322
rect 537294 711002 537326 711238
rect 537562 711002 537646 711238
rect 537882 711002 537914 711238
rect 537294 682954 537914 711002
rect 537294 682718 537326 682954
rect 537562 682718 537646 682954
rect 537882 682718 537914 682954
rect 537294 682634 537914 682718
rect 537294 682398 537326 682634
rect 537562 682398 537646 682634
rect 537882 682398 537914 682634
rect 537294 646954 537914 682398
rect 537294 646718 537326 646954
rect 537562 646718 537646 646954
rect 537882 646718 537914 646954
rect 537294 646634 537914 646718
rect 537294 646398 537326 646634
rect 537562 646398 537646 646634
rect 537882 646398 537914 646634
rect 537294 610954 537914 646398
rect 537294 610718 537326 610954
rect 537562 610718 537646 610954
rect 537882 610718 537914 610954
rect 537294 610634 537914 610718
rect 537294 610398 537326 610634
rect 537562 610398 537646 610634
rect 537882 610398 537914 610634
rect 537294 574954 537914 610398
rect 537294 574718 537326 574954
rect 537562 574718 537646 574954
rect 537882 574718 537914 574954
rect 537294 574634 537914 574718
rect 537294 574398 537326 574634
rect 537562 574398 537646 574634
rect 537882 574398 537914 574634
rect 537294 538954 537914 574398
rect 537294 538718 537326 538954
rect 537562 538718 537646 538954
rect 537882 538718 537914 538954
rect 537294 538634 537914 538718
rect 537294 538398 537326 538634
rect 537562 538398 537646 538634
rect 537882 538398 537914 538634
rect 537294 502954 537914 538398
rect 537294 502718 537326 502954
rect 537562 502718 537646 502954
rect 537882 502718 537914 502954
rect 537294 502634 537914 502718
rect 537294 502398 537326 502634
rect 537562 502398 537646 502634
rect 537882 502398 537914 502634
rect 537294 466954 537914 502398
rect 537294 466718 537326 466954
rect 537562 466718 537646 466954
rect 537882 466718 537914 466954
rect 537294 466634 537914 466718
rect 537294 466398 537326 466634
rect 537562 466398 537646 466634
rect 537882 466398 537914 466634
rect 537294 430954 537914 466398
rect 537294 430718 537326 430954
rect 537562 430718 537646 430954
rect 537882 430718 537914 430954
rect 537294 430634 537914 430718
rect 537294 430398 537326 430634
rect 537562 430398 537646 430634
rect 537882 430398 537914 430634
rect 537294 394954 537914 430398
rect 537294 394718 537326 394954
rect 537562 394718 537646 394954
rect 537882 394718 537914 394954
rect 537294 394634 537914 394718
rect 537294 394398 537326 394634
rect 537562 394398 537646 394634
rect 537882 394398 537914 394634
rect 537294 358954 537914 394398
rect 537294 358718 537326 358954
rect 537562 358718 537646 358954
rect 537882 358718 537914 358954
rect 537294 358634 537914 358718
rect 537294 358398 537326 358634
rect 537562 358398 537646 358634
rect 537882 358398 537914 358634
rect 537294 322954 537914 358398
rect 537294 322718 537326 322954
rect 537562 322718 537646 322954
rect 537882 322718 537914 322954
rect 537294 322634 537914 322718
rect 537294 322398 537326 322634
rect 537562 322398 537646 322634
rect 537882 322398 537914 322634
rect 537294 286954 537914 322398
rect 537294 286718 537326 286954
rect 537562 286718 537646 286954
rect 537882 286718 537914 286954
rect 537294 286634 537914 286718
rect 537294 286398 537326 286634
rect 537562 286398 537646 286634
rect 537882 286398 537914 286634
rect 537294 250954 537914 286398
rect 537294 250718 537326 250954
rect 537562 250718 537646 250954
rect 537882 250718 537914 250954
rect 537294 250634 537914 250718
rect 537294 250398 537326 250634
rect 537562 250398 537646 250634
rect 537882 250398 537914 250634
rect 537294 214954 537914 250398
rect 537294 214718 537326 214954
rect 537562 214718 537646 214954
rect 537882 214718 537914 214954
rect 537294 214634 537914 214718
rect 537294 214398 537326 214634
rect 537562 214398 537646 214634
rect 537882 214398 537914 214634
rect 537294 178954 537914 214398
rect 537294 178718 537326 178954
rect 537562 178718 537646 178954
rect 537882 178718 537914 178954
rect 537294 178634 537914 178718
rect 537294 178398 537326 178634
rect 537562 178398 537646 178634
rect 537882 178398 537914 178634
rect 537294 142954 537914 178398
rect 537294 142718 537326 142954
rect 537562 142718 537646 142954
rect 537882 142718 537914 142954
rect 537294 142634 537914 142718
rect 537294 142398 537326 142634
rect 537562 142398 537646 142634
rect 537882 142398 537914 142634
rect 537294 106954 537914 142398
rect 537294 106718 537326 106954
rect 537562 106718 537646 106954
rect 537882 106718 537914 106954
rect 537294 106634 537914 106718
rect 537294 106398 537326 106634
rect 537562 106398 537646 106634
rect 537882 106398 537914 106634
rect 537294 70954 537914 106398
rect 537294 70718 537326 70954
rect 537562 70718 537646 70954
rect 537882 70718 537914 70954
rect 537294 70634 537914 70718
rect 537294 70398 537326 70634
rect 537562 70398 537646 70634
rect 537882 70398 537914 70634
rect 537294 34954 537914 70398
rect 537294 34718 537326 34954
rect 537562 34718 537646 34954
rect 537882 34718 537914 34954
rect 537294 34634 537914 34718
rect 537294 34398 537326 34634
rect 537562 34398 537646 34634
rect 537882 34398 537914 34634
rect 537294 -7066 537914 34398
rect 537294 -7302 537326 -7066
rect 537562 -7302 537646 -7066
rect 537882 -7302 537914 -7066
rect 537294 -7386 537914 -7302
rect 537294 -7622 537326 -7386
rect 537562 -7622 537646 -7386
rect 537882 -7622 537914 -7386
rect 537294 -7654 537914 -7622
rect 541794 704838 542414 711590
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 687454 542414 704282
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 541794 651454 542414 686898
rect 541794 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 542414 651454
rect 541794 651134 542414 651218
rect 541794 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 542414 651134
rect 541794 615454 542414 650898
rect 541794 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 542414 615454
rect 541794 615134 542414 615218
rect 541794 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 542414 615134
rect 541794 579454 542414 614898
rect 541794 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 542414 579454
rect 541794 579134 542414 579218
rect 541794 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 542414 579134
rect 541794 543454 542414 578898
rect 541794 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 542414 543454
rect 541794 543134 542414 543218
rect 541794 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 542414 543134
rect 541794 507454 542414 542898
rect 541794 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 542414 507454
rect 541794 507134 542414 507218
rect 541794 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 542414 507134
rect 541794 471454 542414 506898
rect 541794 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 542414 471454
rect 541794 471134 542414 471218
rect 541794 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 542414 471134
rect 541794 435454 542414 470898
rect 541794 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 542414 435454
rect 541794 435134 542414 435218
rect 541794 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 542414 435134
rect 541794 399454 542414 434898
rect 541794 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 542414 399454
rect 541794 399134 542414 399218
rect 541794 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 542414 399134
rect 541794 363454 542414 398898
rect 541794 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 542414 363454
rect 541794 363134 542414 363218
rect 541794 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 542414 363134
rect 541794 327454 542414 362898
rect 541794 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 542414 327454
rect 541794 327134 542414 327218
rect 541794 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 542414 327134
rect 541794 291454 542414 326898
rect 541794 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 542414 291454
rect 541794 291134 542414 291218
rect 541794 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 542414 291134
rect 541794 255454 542414 290898
rect 541794 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 542414 255454
rect 541794 255134 542414 255218
rect 541794 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 542414 255134
rect 541794 219454 542414 254898
rect 541794 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 542414 219454
rect 541794 219134 542414 219218
rect 541794 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 542414 219134
rect 541794 183454 542414 218898
rect 541794 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 542414 183454
rect 541794 183134 542414 183218
rect 541794 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 542414 183134
rect 541794 147454 542414 182898
rect 541794 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 542414 147454
rect 541794 147134 542414 147218
rect 541794 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 542414 147134
rect 541794 111454 542414 146898
rect 541794 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 542414 111454
rect 541794 111134 542414 111218
rect 541794 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 542414 111134
rect 541794 75454 542414 110898
rect 541794 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 542414 75454
rect 541794 75134 542414 75218
rect 541794 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 542414 75134
rect 541794 39454 542414 74898
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 541794 3454 542414 38898
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -7654 542414 -902
rect 546294 705798 546914 711590
rect 546294 705562 546326 705798
rect 546562 705562 546646 705798
rect 546882 705562 546914 705798
rect 546294 705478 546914 705562
rect 546294 705242 546326 705478
rect 546562 705242 546646 705478
rect 546882 705242 546914 705478
rect 546294 691954 546914 705242
rect 546294 691718 546326 691954
rect 546562 691718 546646 691954
rect 546882 691718 546914 691954
rect 546294 691634 546914 691718
rect 546294 691398 546326 691634
rect 546562 691398 546646 691634
rect 546882 691398 546914 691634
rect 546294 655954 546914 691398
rect 546294 655718 546326 655954
rect 546562 655718 546646 655954
rect 546882 655718 546914 655954
rect 546294 655634 546914 655718
rect 546294 655398 546326 655634
rect 546562 655398 546646 655634
rect 546882 655398 546914 655634
rect 546294 619954 546914 655398
rect 546294 619718 546326 619954
rect 546562 619718 546646 619954
rect 546882 619718 546914 619954
rect 546294 619634 546914 619718
rect 546294 619398 546326 619634
rect 546562 619398 546646 619634
rect 546882 619398 546914 619634
rect 546294 583954 546914 619398
rect 546294 583718 546326 583954
rect 546562 583718 546646 583954
rect 546882 583718 546914 583954
rect 546294 583634 546914 583718
rect 546294 583398 546326 583634
rect 546562 583398 546646 583634
rect 546882 583398 546914 583634
rect 546294 547954 546914 583398
rect 546294 547718 546326 547954
rect 546562 547718 546646 547954
rect 546882 547718 546914 547954
rect 546294 547634 546914 547718
rect 546294 547398 546326 547634
rect 546562 547398 546646 547634
rect 546882 547398 546914 547634
rect 546294 511954 546914 547398
rect 546294 511718 546326 511954
rect 546562 511718 546646 511954
rect 546882 511718 546914 511954
rect 546294 511634 546914 511718
rect 546294 511398 546326 511634
rect 546562 511398 546646 511634
rect 546882 511398 546914 511634
rect 546294 475954 546914 511398
rect 546294 475718 546326 475954
rect 546562 475718 546646 475954
rect 546882 475718 546914 475954
rect 546294 475634 546914 475718
rect 546294 475398 546326 475634
rect 546562 475398 546646 475634
rect 546882 475398 546914 475634
rect 546294 439954 546914 475398
rect 546294 439718 546326 439954
rect 546562 439718 546646 439954
rect 546882 439718 546914 439954
rect 546294 439634 546914 439718
rect 546294 439398 546326 439634
rect 546562 439398 546646 439634
rect 546882 439398 546914 439634
rect 546294 403954 546914 439398
rect 546294 403718 546326 403954
rect 546562 403718 546646 403954
rect 546882 403718 546914 403954
rect 546294 403634 546914 403718
rect 546294 403398 546326 403634
rect 546562 403398 546646 403634
rect 546882 403398 546914 403634
rect 546294 367954 546914 403398
rect 546294 367718 546326 367954
rect 546562 367718 546646 367954
rect 546882 367718 546914 367954
rect 546294 367634 546914 367718
rect 546294 367398 546326 367634
rect 546562 367398 546646 367634
rect 546882 367398 546914 367634
rect 546294 331954 546914 367398
rect 546294 331718 546326 331954
rect 546562 331718 546646 331954
rect 546882 331718 546914 331954
rect 546294 331634 546914 331718
rect 546294 331398 546326 331634
rect 546562 331398 546646 331634
rect 546882 331398 546914 331634
rect 546294 295954 546914 331398
rect 546294 295718 546326 295954
rect 546562 295718 546646 295954
rect 546882 295718 546914 295954
rect 546294 295634 546914 295718
rect 546294 295398 546326 295634
rect 546562 295398 546646 295634
rect 546882 295398 546914 295634
rect 546294 259954 546914 295398
rect 546294 259718 546326 259954
rect 546562 259718 546646 259954
rect 546882 259718 546914 259954
rect 546294 259634 546914 259718
rect 546294 259398 546326 259634
rect 546562 259398 546646 259634
rect 546882 259398 546914 259634
rect 546294 223954 546914 259398
rect 546294 223718 546326 223954
rect 546562 223718 546646 223954
rect 546882 223718 546914 223954
rect 546294 223634 546914 223718
rect 546294 223398 546326 223634
rect 546562 223398 546646 223634
rect 546882 223398 546914 223634
rect 546294 187954 546914 223398
rect 546294 187718 546326 187954
rect 546562 187718 546646 187954
rect 546882 187718 546914 187954
rect 546294 187634 546914 187718
rect 546294 187398 546326 187634
rect 546562 187398 546646 187634
rect 546882 187398 546914 187634
rect 546294 151954 546914 187398
rect 546294 151718 546326 151954
rect 546562 151718 546646 151954
rect 546882 151718 546914 151954
rect 546294 151634 546914 151718
rect 546294 151398 546326 151634
rect 546562 151398 546646 151634
rect 546882 151398 546914 151634
rect 546294 115954 546914 151398
rect 546294 115718 546326 115954
rect 546562 115718 546646 115954
rect 546882 115718 546914 115954
rect 546294 115634 546914 115718
rect 546294 115398 546326 115634
rect 546562 115398 546646 115634
rect 546882 115398 546914 115634
rect 546294 79954 546914 115398
rect 546294 79718 546326 79954
rect 546562 79718 546646 79954
rect 546882 79718 546914 79954
rect 546294 79634 546914 79718
rect 546294 79398 546326 79634
rect 546562 79398 546646 79634
rect 546882 79398 546914 79634
rect 546294 43954 546914 79398
rect 546294 43718 546326 43954
rect 546562 43718 546646 43954
rect 546882 43718 546914 43954
rect 546294 43634 546914 43718
rect 546294 43398 546326 43634
rect 546562 43398 546646 43634
rect 546882 43398 546914 43634
rect 546294 7954 546914 43398
rect 546294 7718 546326 7954
rect 546562 7718 546646 7954
rect 546882 7718 546914 7954
rect 546294 7634 546914 7718
rect 546294 7398 546326 7634
rect 546562 7398 546646 7634
rect 546882 7398 546914 7634
rect 546294 -1306 546914 7398
rect 546294 -1542 546326 -1306
rect 546562 -1542 546646 -1306
rect 546882 -1542 546914 -1306
rect 546294 -1626 546914 -1542
rect 546294 -1862 546326 -1626
rect 546562 -1862 546646 -1626
rect 546882 -1862 546914 -1626
rect 546294 -7654 546914 -1862
rect 550794 706758 551414 711590
rect 550794 706522 550826 706758
rect 551062 706522 551146 706758
rect 551382 706522 551414 706758
rect 550794 706438 551414 706522
rect 550794 706202 550826 706438
rect 551062 706202 551146 706438
rect 551382 706202 551414 706438
rect 550794 696454 551414 706202
rect 550794 696218 550826 696454
rect 551062 696218 551146 696454
rect 551382 696218 551414 696454
rect 550794 696134 551414 696218
rect 550794 695898 550826 696134
rect 551062 695898 551146 696134
rect 551382 695898 551414 696134
rect 550794 660454 551414 695898
rect 550794 660218 550826 660454
rect 551062 660218 551146 660454
rect 551382 660218 551414 660454
rect 550794 660134 551414 660218
rect 550794 659898 550826 660134
rect 551062 659898 551146 660134
rect 551382 659898 551414 660134
rect 550794 624454 551414 659898
rect 550794 624218 550826 624454
rect 551062 624218 551146 624454
rect 551382 624218 551414 624454
rect 550794 624134 551414 624218
rect 550794 623898 550826 624134
rect 551062 623898 551146 624134
rect 551382 623898 551414 624134
rect 550794 588454 551414 623898
rect 550794 588218 550826 588454
rect 551062 588218 551146 588454
rect 551382 588218 551414 588454
rect 550794 588134 551414 588218
rect 550794 587898 550826 588134
rect 551062 587898 551146 588134
rect 551382 587898 551414 588134
rect 550794 552454 551414 587898
rect 550794 552218 550826 552454
rect 551062 552218 551146 552454
rect 551382 552218 551414 552454
rect 550794 552134 551414 552218
rect 550794 551898 550826 552134
rect 551062 551898 551146 552134
rect 551382 551898 551414 552134
rect 550794 516454 551414 551898
rect 550794 516218 550826 516454
rect 551062 516218 551146 516454
rect 551382 516218 551414 516454
rect 550794 516134 551414 516218
rect 550794 515898 550826 516134
rect 551062 515898 551146 516134
rect 551382 515898 551414 516134
rect 550794 480454 551414 515898
rect 550794 480218 550826 480454
rect 551062 480218 551146 480454
rect 551382 480218 551414 480454
rect 550794 480134 551414 480218
rect 550794 479898 550826 480134
rect 551062 479898 551146 480134
rect 551382 479898 551414 480134
rect 550794 444454 551414 479898
rect 550794 444218 550826 444454
rect 551062 444218 551146 444454
rect 551382 444218 551414 444454
rect 550794 444134 551414 444218
rect 550794 443898 550826 444134
rect 551062 443898 551146 444134
rect 551382 443898 551414 444134
rect 550794 408454 551414 443898
rect 550794 408218 550826 408454
rect 551062 408218 551146 408454
rect 551382 408218 551414 408454
rect 550794 408134 551414 408218
rect 550794 407898 550826 408134
rect 551062 407898 551146 408134
rect 551382 407898 551414 408134
rect 550794 372454 551414 407898
rect 550794 372218 550826 372454
rect 551062 372218 551146 372454
rect 551382 372218 551414 372454
rect 550794 372134 551414 372218
rect 550794 371898 550826 372134
rect 551062 371898 551146 372134
rect 551382 371898 551414 372134
rect 550794 336454 551414 371898
rect 550794 336218 550826 336454
rect 551062 336218 551146 336454
rect 551382 336218 551414 336454
rect 550794 336134 551414 336218
rect 550794 335898 550826 336134
rect 551062 335898 551146 336134
rect 551382 335898 551414 336134
rect 550794 300454 551414 335898
rect 550794 300218 550826 300454
rect 551062 300218 551146 300454
rect 551382 300218 551414 300454
rect 550794 300134 551414 300218
rect 550794 299898 550826 300134
rect 551062 299898 551146 300134
rect 551382 299898 551414 300134
rect 550794 264454 551414 299898
rect 550794 264218 550826 264454
rect 551062 264218 551146 264454
rect 551382 264218 551414 264454
rect 550794 264134 551414 264218
rect 550794 263898 550826 264134
rect 551062 263898 551146 264134
rect 551382 263898 551414 264134
rect 550794 228454 551414 263898
rect 550794 228218 550826 228454
rect 551062 228218 551146 228454
rect 551382 228218 551414 228454
rect 550794 228134 551414 228218
rect 550794 227898 550826 228134
rect 551062 227898 551146 228134
rect 551382 227898 551414 228134
rect 550794 192454 551414 227898
rect 550794 192218 550826 192454
rect 551062 192218 551146 192454
rect 551382 192218 551414 192454
rect 550794 192134 551414 192218
rect 550794 191898 550826 192134
rect 551062 191898 551146 192134
rect 551382 191898 551414 192134
rect 550794 156454 551414 191898
rect 550794 156218 550826 156454
rect 551062 156218 551146 156454
rect 551382 156218 551414 156454
rect 550794 156134 551414 156218
rect 550794 155898 550826 156134
rect 551062 155898 551146 156134
rect 551382 155898 551414 156134
rect 550794 120454 551414 155898
rect 550794 120218 550826 120454
rect 551062 120218 551146 120454
rect 551382 120218 551414 120454
rect 550794 120134 551414 120218
rect 550794 119898 550826 120134
rect 551062 119898 551146 120134
rect 551382 119898 551414 120134
rect 550794 84454 551414 119898
rect 550794 84218 550826 84454
rect 551062 84218 551146 84454
rect 551382 84218 551414 84454
rect 550794 84134 551414 84218
rect 550794 83898 550826 84134
rect 551062 83898 551146 84134
rect 551382 83898 551414 84134
rect 550794 48454 551414 83898
rect 550794 48218 550826 48454
rect 551062 48218 551146 48454
rect 551382 48218 551414 48454
rect 550794 48134 551414 48218
rect 550794 47898 550826 48134
rect 551062 47898 551146 48134
rect 551382 47898 551414 48134
rect 550794 12454 551414 47898
rect 550794 12218 550826 12454
rect 551062 12218 551146 12454
rect 551382 12218 551414 12454
rect 550794 12134 551414 12218
rect 550794 11898 550826 12134
rect 551062 11898 551146 12134
rect 551382 11898 551414 12134
rect 550794 -2266 551414 11898
rect 550794 -2502 550826 -2266
rect 551062 -2502 551146 -2266
rect 551382 -2502 551414 -2266
rect 550794 -2586 551414 -2502
rect 550794 -2822 550826 -2586
rect 551062 -2822 551146 -2586
rect 551382 -2822 551414 -2586
rect 550794 -7654 551414 -2822
rect 555294 707718 555914 711590
rect 555294 707482 555326 707718
rect 555562 707482 555646 707718
rect 555882 707482 555914 707718
rect 555294 707398 555914 707482
rect 555294 707162 555326 707398
rect 555562 707162 555646 707398
rect 555882 707162 555914 707398
rect 555294 700954 555914 707162
rect 555294 700718 555326 700954
rect 555562 700718 555646 700954
rect 555882 700718 555914 700954
rect 555294 700634 555914 700718
rect 555294 700398 555326 700634
rect 555562 700398 555646 700634
rect 555882 700398 555914 700634
rect 555294 664954 555914 700398
rect 555294 664718 555326 664954
rect 555562 664718 555646 664954
rect 555882 664718 555914 664954
rect 555294 664634 555914 664718
rect 555294 664398 555326 664634
rect 555562 664398 555646 664634
rect 555882 664398 555914 664634
rect 555294 628954 555914 664398
rect 555294 628718 555326 628954
rect 555562 628718 555646 628954
rect 555882 628718 555914 628954
rect 555294 628634 555914 628718
rect 555294 628398 555326 628634
rect 555562 628398 555646 628634
rect 555882 628398 555914 628634
rect 555294 592954 555914 628398
rect 555294 592718 555326 592954
rect 555562 592718 555646 592954
rect 555882 592718 555914 592954
rect 555294 592634 555914 592718
rect 555294 592398 555326 592634
rect 555562 592398 555646 592634
rect 555882 592398 555914 592634
rect 555294 556954 555914 592398
rect 555294 556718 555326 556954
rect 555562 556718 555646 556954
rect 555882 556718 555914 556954
rect 555294 556634 555914 556718
rect 555294 556398 555326 556634
rect 555562 556398 555646 556634
rect 555882 556398 555914 556634
rect 555294 520954 555914 556398
rect 555294 520718 555326 520954
rect 555562 520718 555646 520954
rect 555882 520718 555914 520954
rect 555294 520634 555914 520718
rect 555294 520398 555326 520634
rect 555562 520398 555646 520634
rect 555882 520398 555914 520634
rect 555294 484954 555914 520398
rect 555294 484718 555326 484954
rect 555562 484718 555646 484954
rect 555882 484718 555914 484954
rect 555294 484634 555914 484718
rect 555294 484398 555326 484634
rect 555562 484398 555646 484634
rect 555882 484398 555914 484634
rect 555294 448954 555914 484398
rect 555294 448718 555326 448954
rect 555562 448718 555646 448954
rect 555882 448718 555914 448954
rect 555294 448634 555914 448718
rect 555294 448398 555326 448634
rect 555562 448398 555646 448634
rect 555882 448398 555914 448634
rect 555294 412954 555914 448398
rect 555294 412718 555326 412954
rect 555562 412718 555646 412954
rect 555882 412718 555914 412954
rect 555294 412634 555914 412718
rect 555294 412398 555326 412634
rect 555562 412398 555646 412634
rect 555882 412398 555914 412634
rect 555294 376954 555914 412398
rect 555294 376718 555326 376954
rect 555562 376718 555646 376954
rect 555882 376718 555914 376954
rect 555294 376634 555914 376718
rect 555294 376398 555326 376634
rect 555562 376398 555646 376634
rect 555882 376398 555914 376634
rect 555294 340954 555914 376398
rect 555294 340718 555326 340954
rect 555562 340718 555646 340954
rect 555882 340718 555914 340954
rect 555294 340634 555914 340718
rect 555294 340398 555326 340634
rect 555562 340398 555646 340634
rect 555882 340398 555914 340634
rect 555294 304954 555914 340398
rect 555294 304718 555326 304954
rect 555562 304718 555646 304954
rect 555882 304718 555914 304954
rect 555294 304634 555914 304718
rect 555294 304398 555326 304634
rect 555562 304398 555646 304634
rect 555882 304398 555914 304634
rect 555294 268954 555914 304398
rect 555294 268718 555326 268954
rect 555562 268718 555646 268954
rect 555882 268718 555914 268954
rect 555294 268634 555914 268718
rect 555294 268398 555326 268634
rect 555562 268398 555646 268634
rect 555882 268398 555914 268634
rect 555294 232954 555914 268398
rect 555294 232718 555326 232954
rect 555562 232718 555646 232954
rect 555882 232718 555914 232954
rect 555294 232634 555914 232718
rect 555294 232398 555326 232634
rect 555562 232398 555646 232634
rect 555882 232398 555914 232634
rect 555294 196954 555914 232398
rect 555294 196718 555326 196954
rect 555562 196718 555646 196954
rect 555882 196718 555914 196954
rect 555294 196634 555914 196718
rect 555294 196398 555326 196634
rect 555562 196398 555646 196634
rect 555882 196398 555914 196634
rect 555294 160954 555914 196398
rect 555294 160718 555326 160954
rect 555562 160718 555646 160954
rect 555882 160718 555914 160954
rect 555294 160634 555914 160718
rect 555294 160398 555326 160634
rect 555562 160398 555646 160634
rect 555882 160398 555914 160634
rect 555294 124954 555914 160398
rect 555294 124718 555326 124954
rect 555562 124718 555646 124954
rect 555882 124718 555914 124954
rect 555294 124634 555914 124718
rect 555294 124398 555326 124634
rect 555562 124398 555646 124634
rect 555882 124398 555914 124634
rect 555294 88954 555914 124398
rect 555294 88718 555326 88954
rect 555562 88718 555646 88954
rect 555882 88718 555914 88954
rect 555294 88634 555914 88718
rect 555294 88398 555326 88634
rect 555562 88398 555646 88634
rect 555882 88398 555914 88634
rect 555294 52954 555914 88398
rect 555294 52718 555326 52954
rect 555562 52718 555646 52954
rect 555882 52718 555914 52954
rect 555294 52634 555914 52718
rect 555294 52398 555326 52634
rect 555562 52398 555646 52634
rect 555882 52398 555914 52634
rect 555294 16954 555914 52398
rect 555294 16718 555326 16954
rect 555562 16718 555646 16954
rect 555882 16718 555914 16954
rect 555294 16634 555914 16718
rect 555294 16398 555326 16634
rect 555562 16398 555646 16634
rect 555882 16398 555914 16634
rect 555294 -3226 555914 16398
rect 555294 -3462 555326 -3226
rect 555562 -3462 555646 -3226
rect 555882 -3462 555914 -3226
rect 555294 -3546 555914 -3462
rect 555294 -3782 555326 -3546
rect 555562 -3782 555646 -3546
rect 555882 -3782 555914 -3546
rect 555294 -7654 555914 -3782
rect 559794 708678 560414 711590
rect 559794 708442 559826 708678
rect 560062 708442 560146 708678
rect 560382 708442 560414 708678
rect 559794 708358 560414 708442
rect 559794 708122 559826 708358
rect 560062 708122 560146 708358
rect 560382 708122 560414 708358
rect 559794 669454 560414 708122
rect 559794 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 560414 669454
rect 559794 669134 560414 669218
rect 559794 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 560414 669134
rect 559794 633454 560414 668898
rect 559794 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 560414 633454
rect 559794 633134 560414 633218
rect 559794 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 560414 633134
rect 559794 597454 560414 632898
rect 559794 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 560414 597454
rect 559794 597134 560414 597218
rect 559794 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 560414 597134
rect 559794 561454 560414 596898
rect 559794 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 560414 561454
rect 559794 561134 560414 561218
rect 559794 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 560414 561134
rect 559794 525454 560414 560898
rect 559794 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 560414 525454
rect 559794 525134 560414 525218
rect 559794 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 560414 525134
rect 559794 489454 560414 524898
rect 559794 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 560414 489454
rect 559794 489134 560414 489218
rect 559794 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 560414 489134
rect 559794 453454 560414 488898
rect 559794 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 560414 453454
rect 559794 453134 560414 453218
rect 559794 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 560414 453134
rect 559794 417454 560414 452898
rect 559794 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 560414 417454
rect 559794 417134 560414 417218
rect 559794 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 560414 417134
rect 559794 381454 560414 416898
rect 559794 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 560414 381454
rect 559794 381134 560414 381218
rect 559794 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 560414 381134
rect 559794 345454 560414 380898
rect 559794 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 560414 345454
rect 559794 345134 560414 345218
rect 559794 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 560414 345134
rect 559794 309454 560414 344898
rect 559794 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 560414 309454
rect 559794 309134 560414 309218
rect 559794 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 560414 309134
rect 559794 273454 560414 308898
rect 559794 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 560414 273454
rect 559794 273134 560414 273218
rect 559794 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 560414 273134
rect 559794 237454 560414 272898
rect 559794 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 560414 237454
rect 559794 237134 560414 237218
rect 559794 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 560414 237134
rect 559794 201454 560414 236898
rect 559794 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 560414 201454
rect 559794 201134 560414 201218
rect 559794 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 560414 201134
rect 559794 165454 560414 200898
rect 559794 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 560414 165454
rect 559794 165134 560414 165218
rect 559794 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 560414 165134
rect 559794 129454 560414 164898
rect 559794 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 560414 129454
rect 559794 129134 560414 129218
rect 559794 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 560414 129134
rect 559794 93454 560414 128898
rect 559794 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 560414 93454
rect 559794 93134 560414 93218
rect 559794 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 560414 93134
rect 559794 57454 560414 92898
rect 559794 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 560414 57454
rect 559794 57134 560414 57218
rect 559794 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 560414 57134
rect 559794 21454 560414 56898
rect 559794 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 560414 21454
rect 559794 21134 560414 21218
rect 559794 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 560414 21134
rect 559794 -4186 560414 20898
rect 559794 -4422 559826 -4186
rect 560062 -4422 560146 -4186
rect 560382 -4422 560414 -4186
rect 559794 -4506 560414 -4422
rect 559794 -4742 559826 -4506
rect 560062 -4742 560146 -4506
rect 560382 -4742 560414 -4506
rect 559794 -7654 560414 -4742
rect 564294 709638 564914 711590
rect 564294 709402 564326 709638
rect 564562 709402 564646 709638
rect 564882 709402 564914 709638
rect 564294 709318 564914 709402
rect 564294 709082 564326 709318
rect 564562 709082 564646 709318
rect 564882 709082 564914 709318
rect 564294 673954 564914 709082
rect 564294 673718 564326 673954
rect 564562 673718 564646 673954
rect 564882 673718 564914 673954
rect 564294 673634 564914 673718
rect 564294 673398 564326 673634
rect 564562 673398 564646 673634
rect 564882 673398 564914 673634
rect 564294 637954 564914 673398
rect 564294 637718 564326 637954
rect 564562 637718 564646 637954
rect 564882 637718 564914 637954
rect 564294 637634 564914 637718
rect 564294 637398 564326 637634
rect 564562 637398 564646 637634
rect 564882 637398 564914 637634
rect 564294 601954 564914 637398
rect 564294 601718 564326 601954
rect 564562 601718 564646 601954
rect 564882 601718 564914 601954
rect 564294 601634 564914 601718
rect 564294 601398 564326 601634
rect 564562 601398 564646 601634
rect 564882 601398 564914 601634
rect 564294 565954 564914 601398
rect 564294 565718 564326 565954
rect 564562 565718 564646 565954
rect 564882 565718 564914 565954
rect 564294 565634 564914 565718
rect 564294 565398 564326 565634
rect 564562 565398 564646 565634
rect 564882 565398 564914 565634
rect 564294 529954 564914 565398
rect 564294 529718 564326 529954
rect 564562 529718 564646 529954
rect 564882 529718 564914 529954
rect 564294 529634 564914 529718
rect 564294 529398 564326 529634
rect 564562 529398 564646 529634
rect 564882 529398 564914 529634
rect 564294 493954 564914 529398
rect 564294 493718 564326 493954
rect 564562 493718 564646 493954
rect 564882 493718 564914 493954
rect 564294 493634 564914 493718
rect 564294 493398 564326 493634
rect 564562 493398 564646 493634
rect 564882 493398 564914 493634
rect 564294 457954 564914 493398
rect 564294 457718 564326 457954
rect 564562 457718 564646 457954
rect 564882 457718 564914 457954
rect 564294 457634 564914 457718
rect 564294 457398 564326 457634
rect 564562 457398 564646 457634
rect 564882 457398 564914 457634
rect 564294 421954 564914 457398
rect 564294 421718 564326 421954
rect 564562 421718 564646 421954
rect 564882 421718 564914 421954
rect 564294 421634 564914 421718
rect 564294 421398 564326 421634
rect 564562 421398 564646 421634
rect 564882 421398 564914 421634
rect 564294 385954 564914 421398
rect 564294 385718 564326 385954
rect 564562 385718 564646 385954
rect 564882 385718 564914 385954
rect 564294 385634 564914 385718
rect 564294 385398 564326 385634
rect 564562 385398 564646 385634
rect 564882 385398 564914 385634
rect 564294 349954 564914 385398
rect 564294 349718 564326 349954
rect 564562 349718 564646 349954
rect 564882 349718 564914 349954
rect 564294 349634 564914 349718
rect 564294 349398 564326 349634
rect 564562 349398 564646 349634
rect 564882 349398 564914 349634
rect 564294 313954 564914 349398
rect 564294 313718 564326 313954
rect 564562 313718 564646 313954
rect 564882 313718 564914 313954
rect 564294 313634 564914 313718
rect 564294 313398 564326 313634
rect 564562 313398 564646 313634
rect 564882 313398 564914 313634
rect 564294 277954 564914 313398
rect 564294 277718 564326 277954
rect 564562 277718 564646 277954
rect 564882 277718 564914 277954
rect 564294 277634 564914 277718
rect 564294 277398 564326 277634
rect 564562 277398 564646 277634
rect 564882 277398 564914 277634
rect 564294 241954 564914 277398
rect 564294 241718 564326 241954
rect 564562 241718 564646 241954
rect 564882 241718 564914 241954
rect 564294 241634 564914 241718
rect 564294 241398 564326 241634
rect 564562 241398 564646 241634
rect 564882 241398 564914 241634
rect 564294 205954 564914 241398
rect 564294 205718 564326 205954
rect 564562 205718 564646 205954
rect 564882 205718 564914 205954
rect 564294 205634 564914 205718
rect 564294 205398 564326 205634
rect 564562 205398 564646 205634
rect 564882 205398 564914 205634
rect 564294 169954 564914 205398
rect 564294 169718 564326 169954
rect 564562 169718 564646 169954
rect 564882 169718 564914 169954
rect 564294 169634 564914 169718
rect 564294 169398 564326 169634
rect 564562 169398 564646 169634
rect 564882 169398 564914 169634
rect 564294 133954 564914 169398
rect 564294 133718 564326 133954
rect 564562 133718 564646 133954
rect 564882 133718 564914 133954
rect 564294 133634 564914 133718
rect 564294 133398 564326 133634
rect 564562 133398 564646 133634
rect 564882 133398 564914 133634
rect 564294 97954 564914 133398
rect 564294 97718 564326 97954
rect 564562 97718 564646 97954
rect 564882 97718 564914 97954
rect 564294 97634 564914 97718
rect 564294 97398 564326 97634
rect 564562 97398 564646 97634
rect 564882 97398 564914 97634
rect 564294 61954 564914 97398
rect 564294 61718 564326 61954
rect 564562 61718 564646 61954
rect 564882 61718 564914 61954
rect 564294 61634 564914 61718
rect 564294 61398 564326 61634
rect 564562 61398 564646 61634
rect 564882 61398 564914 61634
rect 564294 25954 564914 61398
rect 564294 25718 564326 25954
rect 564562 25718 564646 25954
rect 564882 25718 564914 25954
rect 564294 25634 564914 25718
rect 564294 25398 564326 25634
rect 564562 25398 564646 25634
rect 564882 25398 564914 25634
rect 564294 -5146 564914 25398
rect 564294 -5382 564326 -5146
rect 564562 -5382 564646 -5146
rect 564882 -5382 564914 -5146
rect 564294 -5466 564914 -5382
rect 564294 -5702 564326 -5466
rect 564562 -5702 564646 -5466
rect 564882 -5702 564914 -5466
rect 564294 -7654 564914 -5702
rect 568794 710598 569414 711590
rect 568794 710362 568826 710598
rect 569062 710362 569146 710598
rect 569382 710362 569414 710598
rect 568794 710278 569414 710362
rect 568794 710042 568826 710278
rect 569062 710042 569146 710278
rect 569382 710042 569414 710278
rect 568794 678454 569414 710042
rect 568794 678218 568826 678454
rect 569062 678218 569146 678454
rect 569382 678218 569414 678454
rect 568794 678134 569414 678218
rect 568794 677898 568826 678134
rect 569062 677898 569146 678134
rect 569382 677898 569414 678134
rect 568794 642454 569414 677898
rect 568794 642218 568826 642454
rect 569062 642218 569146 642454
rect 569382 642218 569414 642454
rect 568794 642134 569414 642218
rect 568794 641898 568826 642134
rect 569062 641898 569146 642134
rect 569382 641898 569414 642134
rect 568794 606454 569414 641898
rect 568794 606218 568826 606454
rect 569062 606218 569146 606454
rect 569382 606218 569414 606454
rect 568794 606134 569414 606218
rect 568794 605898 568826 606134
rect 569062 605898 569146 606134
rect 569382 605898 569414 606134
rect 568794 570454 569414 605898
rect 568794 570218 568826 570454
rect 569062 570218 569146 570454
rect 569382 570218 569414 570454
rect 568794 570134 569414 570218
rect 568794 569898 568826 570134
rect 569062 569898 569146 570134
rect 569382 569898 569414 570134
rect 568794 534454 569414 569898
rect 568794 534218 568826 534454
rect 569062 534218 569146 534454
rect 569382 534218 569414 534454
rect 568794 534134 569414 534218
rect 568794 533898 568826 534134
rect 569062 533898 569146 534134
rect 569382 533898 569414 534134
rect 568794 498454 569414 533898
rect 568794 498218 568826 498454
rect 569062 498218 569146 498454
rect 569382 498218 569414 498454
rect 568794 498134 569414 498218
rect 568794 497898 568826 498134
rect 569062 497898 569146 498134
rect 569382 497898 569414 498134
rect 568794 462454 569414 497898
rect 568794 462218 568826 462454
rect 569062 462218 569146 462454
rect 569382 462218 569414 462454
rect 568794 462134 569414 462218
rect 568794 461898 568826 462134
rect 569062 461898 569146 462134
rect 569382 461898 569414 462134
rect 568794 426454 569414 461898
rect 568794 426218 568826 426454
rect 569062 426218 569146 426454
rect 569382 426218 569414 426454
rect 568794 426134 569414 426218
rect 568794 425898 568826 426134
rect 569062 425898 569146 426134
rect 569382 425898 569414 426134
rect 568794 390454 569414 425898
rect 568794 390218 568826 390454
rect 569062 390218 569146 390454
rect 569382 390218 569414 390454
rect 568794 390134 569414 390218
rect 568794 389898 568826 390134
rect 569062 389898 569146 390134
rect 569382 389898 569414 390134
rect 568794 354454 569414 389898
rect 568794 354218 568826 354454
rect 569062 354218 569146 354454
rect 569382 354218 569414 354454
rect 568794 354134 569414 354218
rect 568794 353898 568826 354134
rect 569062 353898 569146 354134
rect 569382 353898 569414 354134
rect 568794 318454 569414 353898
rect 568794 318218 568826 318454
rect 569062 318218 569146 318454
rect 569382 318218 569414 318454
rect 568794 318134 569414 318218
rect 568794 317898 568826 318134
rect 569062 317898 569146 318134
rect 569382 317898 569414 318134
rect 568794 282454 569414 317898
rect 568794 282218 568826 282454
rect 569062 282218 569146 282454
rect 569382 282218 569414 282454
rect 568794 282134 569414 282218
rect 568794 281898 568826 282134
rect 569062 281898 569146 282134
rect 569382 281898 569414 282134
rect 568794 246454 569414 281898
rect 568794 246218 568826 246454
rect 569062 246218 569146 246454
rect 569382 246218 569414 246454
rect 568794 246134 569414 246218
rect 568794 245898 568826 246134
rect 569062 245898 569146 246134
rect 569382 245898 569414 246134
rect 568794 210454 569414 245898
rect 568794 210218 568826 210454
rect 569062 210218 569146 210454
rect 569382 210218 569414 210454
rect 568794 210134 569414 210218
rect 568794 209898 568826 210134
rect 569062 209898 569146 210134
rect 569382 209898 569414 210134
rect 568794 174454 569414 209898
rect 568794 174218 568826 174454
rect 569062 174218 569146 174454
rect 569382 174218 569414 174454
rect 568794 174134 569414 174218
rect 568794 173898 568826 174134
rect 569062 173898 569146 174134
rect 569382 173898 569414 174134
rect 568794 138454 569414 173898
rect 568794 138218 568826 138454
rect 569062 138218 569146 138454
rect 569382 138218 569414 138454
rect 568794 138134 569414 138218
rect 568794 137898 568826 138134
rect 569062 137898 569146 138134
rect 569382 137898 569414 138134
rect 568794 102454 569414 137898
rect 568794 102218 568826 102454
rect 569062 102218 569146 102454
rect 569382 102218 569414 102454
rect 568794 102134 569414 102218
rect 568794 101898 568826 102134
rect 569062 101898 569146 102134
rect 569382 101898 569414 102134
rect 568794 66454 569414 101898
rect 568794 66218 568826 66454
rect 569062 66218 569146 66454
rect 569382 66218 569414 66454
rect 568794 66134 569414 66218
rect 568794 65898 568826 66134
rect 569062 65898 569146 66134
rect 569382 65898 569414 66134
rect 568794 30454 569414 65898
rect 568794 30218 568826 30454
rect 569062 30218 569146 30454
rect 569382 30218 569414 30454
rect 568794 30134 569414 30218
rect 568794 29898 568826 30134
rect 569062 29898 569146 30134
rect 569382 29898 569414 30134
rect 568794 -6106 569414 29898
rect 568794 -6342 568826 -6106
rect 569062 -6342 569146 -6106
rect 569382 -6342 569414 -6106
rect 568794 -6426 569414 -6342
rect 568794 -6662 568826 -6426
rect 569062 -6662 569146 -6426
rect 569382 -6662 569414 -6426
rect 568794 -7654 569414 -6662
rect 573294 711558 573914 711590
rect 573294 711322 573326 711558
rect 573562 711322 573646 711558
rect 573882 711322 573914 711558
rect 573294 711238 573914 711322
rect 573294 711002 573326 711238
rect 573562 711002 573646 711238
rect 573882 711002 573914 711238
rect 573294 682954 573914 711002
rect 573294 682718 573326 682954
rect 573562 682718 573646 682954
rect 573882 682718 573914 682954
rect 573294 682634 573914 682718
rect 573294 682398 573326 682634
rect 573562 682398 573646 682634
rect 573882 682398 573914 682634
rect 573294 646954 573914 682398
rect 573294 646718 573326 646954
rect 573562 646718 573646 646954
rect 573882 646718 573914 646954
rect 573294 646634 573914 646718
rect 573294 646398 573326 646634
rect 573562 646398 573646 646634
rect 573882 646398 573914 646634
rect 573294 610954 573914 646398
rect 573294 610718 573326 610954
rect 573562 610718 573646 610954
rect 573882 610718 573914 610954
rect 573294 610634 573914 610718
rect 573294 610398 573326 610634
rect 573562 610398 573646 610634
rect 573882 610398 573914 610634
rect 573294 574954 573914 610398
rect 573294 574718 573326 574954
rect 573562 574718 573646 574954
rect 573882 574718 573914 574954
rect 573294 574634 573914 574718
rect 573294 574398 573326 574634
rect 573562 574398 573646 574634
rect 573882 574398 573914 574634
rect 573294 538954 573914 574398
rect 573294 538718 573326 538954
rect 573562 538718 573646 538954
rect 573882 538718 573914 538954
rect 573294 538634 573914 538718
rect 573294 538398 573326 538634
rect 573562 538398 573646 538634
rect 573882 538398 573914 538634
rect 573294 502954 573914 538398
rect 573294 502718 573326 502954
rect 573562 502718 573646 502954
rect 573882 502718 573914 502954
rect 573294 502634 573914 502718
rect 573294 502398 573326 502634
rect 573562 502398 573646 502634
rect 573882 502398 573914 502634
rect 573294 466954 573914 502398
rect 573294 466718 573326 466954
rect 573562 466718 573646 466954
rect 573882 466718 573914 466954
rect 573294 466634 573914 466718
rect 573294 466398 573326 466634
rect 573562 466398 573646 466634
rect 573882 466398 573914 466634
rect 573294 430954 573914 466398
rect 573294 430718 573326 430954
rect 573562 430718 573646 430954
rect 573882 430718 573914 430954
rect 573294 430634 573914 430718
rect 573294 430398 573326 430634
rect 573562 430398 573646 430634
rect 573882 430398 573914 430634
rect 573294 394954 573914 430398
rect 573294 394718 573326 394954
rect 573562 394718 573646 394954
rect 573882 394718 573914 394954
rect 573294 394634 573914 394718
rect 573294 394398 573326 394634
rect 573562 394398 573646 394634
rect 573882 394398 573914 394634
rect 573294 358954 573914 394398
rect 573294 358718 573326 358954
rect 573562 358718 573646 358954
rect 573882 358718 573914 358954
rect 573294 358634 573914 358718
rect 573294 358398 573326 358634
rect 573562 358398 573646 358634
rect 573882 358398 573914 358634
rect 573294 322954 573914 358398
rect 573294 322718 573326 322954
rect 573562 322718 573646 322954
rect 573882 322718 573914 322954
rect 573294 322634 573914 322718
rect 573294 322398 573326 322634
rect 573562 322398 573646 322634
rect 573882 322398 573914 322634
rect 573294 286954 573914 322398
rect 573294 286718 573326 286954
rect 573562 286718 573646 286954
rect 573882 286718 573914 286954
rect 573294 286634 573914 286718
rect 573294 286398 573326 286634
rect 573562 286398 573646 286634
rect 573882 286398 573914 286634
rect 573294 250954 573914 286398
rect 573294 250718 573326 250954
rect 573562 250718 573646 250954
rect 573882 250718 573914 250954
rect 573294 250634 573914 250718
rect 573294 250398 573326 250634
rect 573562 250398 573646 250634
rect 573882 250398 573914 250634
rect 573294 214954 573914 250398
rect 573294 214718 573326 214954
rect 573562 214718 573646 214954
rect 573882 214718 573914 214954
rect 573294 214634 573914 214718
rect 573294 214398 573326 214634
rect 573562 214398 573646 214634
rect 573882 214398 573914 214634
rect 573294 178954 573914 214398
rect 573294 178718 573326 178954
rect 573562 178718 573646 178954
rect 573882 178718 573914 178954
rect 573294 178634 573914 178718
rect 573294 178398 573326 178634
rect 573562 178398 573646 178634
rect 573882 178398 573914 178634
rect 573294 142954 573914 178398
rect 573294 142718 573326 142954
rect 573562 142718 573646 142954
rect 573882 142718 573914 142954
rect 573294 142634 573914 142718
rect 573294 142398 573326 142634
rect 573562 142398 573646 142634
rect 573882 142398 573914 142634
rect 573294 106954 573914 142398
rect 573294 106718 573326 106954
rect 573562 106718 573646 106954
rect 573882 106718 573914 106954
rect 573294 106634 573914 106718
rect 573294 106398 573326 106634
rect 573562 106398 573646 106634
rect 573882 106398 573914 106634
rect 573294 70954 573914 106398
rect 573294 70718 573326 70954
rect 573562 70718 573646 70954
rect 573882 70718 573914 70954
rect 573294 70634 573914 70718
rect 573294 70398 573326 70634
rect 573562 70398 573646 70634
rect 573882 70398 573914 70634
rect 573294 34954 573914 70398
rect 573294 34718 573326 34954
rect 573562 34718 573646 34954
rect 573882 34718 573914 34954
rect 573294 34634 573914 34718
rect 573294 34398 573326 34634
rect 573562 34398 573646 34634
rect 573882 34398 573914 34634
rect 573294 -7066 573914 34398
rect 573294 -7302 573326 -7066
rect 573562 -7302 573646 -7066
rect 573882 -7302 573914 -7066
rect 573294 -7386 573914 -7302
rect 573294 -7622 573326 -7386
rect 573562 -7622 573646 -7386
rect 573882 -7622 573914 -7386
rect 573294 -7654 573914 -7622
rect 577794 704838 578414 711590
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 582294 705798 582914 711590
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 582294 705562 582326 705798
rect 582562 705562 582646 705798
rect 582882 705562 582914 705798
rect 582294 705478 582914 705562
rect 582294 705242 582326 705478
rect 582562 705242 582646 705478
rect 582882 705242 582914 705478
rect 582294 691954 582914 705242
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 582294 691718 582326 691954
rect 582562 691718 582646 691954
rect 582882 691718 582914 691954
rect 582294 691634 582914 691718
rect 582294 691398 582326 691634
rect 582562 691398 582646 691634
rect 582882 691398 582914 691634
rect 582294 655954 582914 691398
rect 582294 655718 582326 655954
rect 582562 655718 582646 655954
rect 582882 655718 582914 655954
rect 582294 655634 582914 655718
rect 582294 655398 582326 655634
rect 582562 655398 582646 655634
rect 582882 655398 582914 655634
rect 582294 619954 582914 655398
rect 582294 619718 582326 619954
rect 582562 619718 582646 619954
rect 582882 619718 582914 619954
rect 582294 619634 582914 619718
rect 582294 619398 582326 619634
rect 582562 619398 582646 619634
rect 582882 619398 582914 619634
rect 582294 583954 582914 619398
rect 582294 583718 582326 583954
rect 582562 583718 582646 583954
rect 582882 583718 582914 583954
rect 582294 583634 582914 583718
rect 582294 583398 582326 583634
rect 582562 583398 582646 583634
rect 582882 583398 582914 583634
rect 582294 547954 582914 583398
rect 582294 547718 582326 547954
rect 582562 547718 582646 547954
rect 582882 547718 582914 547954
rect 582294 547634 582914 547718
rect 582294 547398 582326 547634
rect 582562 547398 582646 547634
rect 582882 547398 582914 547634
rect 582294 511954 582914 547398
rect 582294 511718 582326 511954
rect 582562 511718 582646 511954
rect 582882 511718 582914 511954
rect 582294 511634 582914 511718
rect 582294 511398 582326 511634
rect 582562 511398 582646 511634
rect 582882 511398 582914 511634
rect 582294 475954 582914 511398
rect 582294 475718 582326 475954
rect 582562 475718 582646 475954
rect 582882 475718 582914 475954
rect 582294 475634 582914 475718
rect 582294 475398 582326 475634
rect 582562 475398 582646 475634
rect 582882 475398 582914 475634
rect 582294 439954 582914 475398
rect 582294 439718 582326 439954
rect 582562 439718 582646 439954
rect 582882 439718 582914 439954
rect 582294 439634 582914 439718
rect 582294 439398 582326 439634
rect 582562 439398 582646 439634
rect 582882 439398 582914 439634
rect 582294 403954 582914 439398
rect 582294 403718 582326 403954
rect 582562 403718 582646 403954
rect 582882 403718 582914 403954
rect 582294 403634 582914 403718
rect 582294 403398 582326 403634
rect 582562 403398 582646 403634
rect 582882 403398 582914 403634
rect 580211 381580 580277 381581
rect 580211 381516 580212 381580
rect 580276 381516 580277 381580
rect 580211 381515 580277 381516
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 580214 59669 580274 381515
rect 582294 367954 582914 403398
rect 582294 367718 582326 367954
rect 582562 367718 582646 367954
rect 582882 367718 582914 367954
rect 582294 367634 582914 367718
rect 582294 367398 582326 367634
rect 582562 367398 582646 367634
rect 582882 367398 582914 367634
rect 582294 331954 582914 367398
rect 582294 331718 582326 331954
rect 582562 331718 582646 331954
rect 582882 331718 582914 331954
rect 582294 331634 582914 331718
rect 582294 331398 582326 331634
rect 582562 331398 582646 331634
rect 582882 331398 582914 331634
rect 582294 295954 582914 331398
rect 582294 295718 582326 295954
rect 582562 295718 582646 295954
rect 582882 295718 582914 295954
rect 582294 295634 582914 295718
rect 582294 295398 582326 295634
rect 582562 295398 582646 295634
rect 582882 295398 582914 295634
rect 582294 259954 582914 295398
rect 582294 259718 582326 259954
rect 582562 259718 582646 259954
rect 582882 259718 582914 259954
rect 582294 259634 582914 259718
rect 582294 259398 582326 259634
rect 582562 259398 582646 259634
rect 582882 259398 582914 259634
rect 582294 223954 582914 259398
rect 582294 223718 582326 223954
rect 582562 223718 582646 223954
rect 582882 223718 582914 223954
rect 582294 223634 582914 223718
rect 582294 223398 582326 223634
rect 582562 223398 582646 223634
rect 582882 223398 582914 223634
rect 582294 187954 582914 223398
rect 582294 187718 582326 187954
rect 582562 187718 582646 187954
rect 582882 187718 582914 187954
rect 582294 187634 582914 187718
rect 582294 187398 582326 187634
rect 582562 187398 582646 187634
rect 582882 187398 582914 187634
rect 582294 151954 582914 187398
rect 582294 151718 582326 151954
rect 582562 151718 582646 151954
rect 582882 151718 582914 151954
rect 582294 151634 582914 151718
rect 582294 151398 582326 151634
rect 582562 151398 582646 151634
rect 582882 151398 582914 151634
rect 582294 115954 582914 151398
rect 582294 115718 582326 115954
rect 582562 115718 582646 115954
rect 582882 115718 582914 115954
rect 582294 115634 582914 115718
rect 582294 115398 582326 115634
rect 582562 115398 582646 115634
rect 582882 115398 582914 115634
rect 582294 79954 582914 115398
rect 582294 79718 582326 79954
rect 582562 79718 582646 79954
rect 582882 79718 582914 79954
rect 582294 79634 582914 79718
rect 582294 79398 582326 79634
rect 582562 79398 582646 79634
rect 582882 79398 582914 79634
rect 580211 59668 580277 59669
rect 580211 59604 580212 59668
rect 580276 59604 580277 59668
rect 580211 59603 580277 59604
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -7654 578414 -902
rect 582294 43954 582914 79398
rect 582294 43718 582326 43954
rect 582562 43718 582646 43954
rect 582882 43718 582914 43954
rect 582294 43634 582914 43718
rect 582294 43398 582326 43634
rect 582562 43398 582646 43634
rect 582882 43398 582914 43634
rect 582294 7954 582914 43398
rect 582294 7718 582326 7954
rect 582562 7718 582646 7954
rect 582882 7718 582914 7954
rect 582294 7634 582914 7718
rect 582294 7398 582326 7634
rect 582562 7398 582646 7634
rect 582882 7398 582914 7634
rect 582294 -1306 582914 7398
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 691954 586890 705242
rect 586270 691718 586302 691954
rect 586538 691718 586622 691954
rect 586858 691718 586890 691954
rect 586270 691634 586890 691718
rect 586270 691398 586302 691634
rect 586538 691398 586622 691634
rect 586858 691398 586890 691634
rect 586270 655954 586890 691398
rect 586270 655718 586302 655954
rect 586538 655718 586622 655954
rect 586858 655718 586890 655954
rect 586270 655634 586890 655718
rect 586270 655398 586302 655634
rect 586538 655398 586622 655634
rect 586858 655398 586890 655634
rect 586270 619954 586890 655398
rect 586270 619718 586302 619954
rect 586538 619718 586622 619954
rect 586858 619718 586890 619954
rect 586270 619634 586890 619718
rect 586270 619398 586302 619634
rect 586538 619398 586622 619634
rect 586858 619398 586890 619634
rect 586270 583954 586890 619398
rect 586270 583718 586302 583954
rect 586538 583718 586622 583954
rect 586858 583718 586890 583954
rect 586270 583634 586890 583718
rect 586270 583398 586302 583634
rect 586538 583398 586622 583634
rect 586858 583398 586890 583634
rect 586270 547954 586890 583398
rect 586270 547718 586302 547954
rect 586538 547718 586622 547954
rect 586858 547718 586890 547954
rect 586270 547634 586890 547718
rect 586270 547398 586302 547634
rect 586538 547398 586622 547634
rect 586858 547398 586890 547634
rect 586270 511954 586890 547398
rect 586270 511718 586302 511954
rect 586538 511718 586622 511954
rect 586858 511718 586890 511954
rect 586270 511634 586890 511718
rect 586270 511398 586302 511634
rect 586538 511398 586622 511634
rect 586858 511398 586890 511634
rect 586270 475954 586890 511398
rect 586270 475718 586302 475954
rect 586538 475718 586622 475954
rect 586858 475718 586890 475954
rect 586270 475634 586890 475718
rect 586270 475398 586302 475634
rect 586538 475398 586622 475634
rect 586858 475398 586890 475634
rect 586270 439954 586890 475398
rect 586270 439718 586302 439954
rect 586538 439718 586622 439954
rect 586858 439718 586890 439954
rect 586270 439634 586890 439718
rect 586270 439398 586302 439634
rect 586538 439398 586622 439634
rect 586858 439398 586890 439634
rect 586270 403954 586890 439398
rect 586270 403718 586302 403954
rect 586538 403718 586622 403954
rect 586858 403718 586890 403954
rect 586270 403634 586890 403718
rect 586270 403398 586302 403634
rect 586538 403398 586622 403634
rect 586858 403398 586890 403634
rect 586270 367954 586890 403398
rect 586270 367718 586302 367954
rect 586538 367718 586622 367954
rect 586858 367718 586890 367954
rect 586270 367634 586890 367718
rect 586270 367398 586302 367634
rect 586538 367398 586622 367634
rect 586858 367398 586890 367634
rect 586270 331954 586890 367398
rect 586270 331718 586302 331954
rect 586538 331718 586622 331954
rect 586858 331718 586890 331954
rect 586270 331634 586890 331718
rect 586270 331398 586302 331634
rect 586538 331398 586622 331634
rect 586858 331398 586890 331634
rect 586270 295954 586890 331398
rect 586270 295718 586302 295954
rect 586538 295718 586622 295954
rect 586858 295718 586890 295954
rect 586270 295634 586890 295718
rect 586270 295398 586302 295634
rect 586538 295398 586622 295634
rect 586858 295398 586890 295634
rect 586270 259954 586890 295398
rect 586270 259718 586302 259954
rect 586538 259718 586622 259954
rect 586858 259718 586890 259954
rect 586270 259634 586890 259718
rect 586270 259398 586302 259634
rect 586538 259398 586622 259634
rect 586858 259398 586890 259634
rect 586270 223954 586890 259398
rect 586270 223718 586302 223954
rect 586538 223718 586622 223954
rect 586858 223718 586890 223954
rect 586270 223634 586890 223718
rect 586270 223398 586302 223634
rect 586538 223398 586622 223634
rect 586858 223398 586890 223634
rect 586270 187954 586890 223398
rect 586270 187718 586302 187954
rect 586538 187718 586622 187954
rect 586858 187718 586890 187954
rect 586270 187634 586890 187718
rect 586270 187398 586302 187634
rect 586538 187398 586622 187634
rect 586858 187398 586890 187634
rect 586270 151954 586890 187398
rect 586270 151718 586302 151954
rect 586538 151718 586622 151954
rect 586858 151718 586890 151954
rect 586270 151634 586890 151718
rect 586270 151398 586302 151634
rect 586538 151398 586622 151634
rect 586858 151398 586890 151634
rect 586270 115954 586890 151398
rect 586270 115718 586302 115954
rect 586538 115718 586622 115954
rect 586858 115718 586890 115954
rect 586270 115634 586890 115718
rect 586270 115398 586302 115634
rect 586538 115398 586622 115634
rect 586858 115398 586890 115634
rect 586270 79954 586890 115398
rect 586270 79718 586302 79954
rect 586538 79718 586622 79954
rect 586858 79718 586890 79954
rect 586270 79634 586890 79718
rect 586270 79398 586302 79634
rect 586538 79398 586622 79634
rect 586858 79398 586890 79634
rect 586270 43954 586890 79398
rect 586270 43718 586302 43954
rect 586538 43718 586622 43954
rect 586858 43718 586890 43954
rect 586270 43634 586890 43718
rect 586270 43398 586302 43634
rect 586538 43398 586622 43634
rect 586858 43398 586890 43634
rect 586270 7954 586890 43398
rect 586270 7718 586302 7954
rect 586538 7718 586622 7954
rect 586858 7718 586890 7954
rect 586270 7634 586890 7718
rect 586270 7398 586302 7634
rect 586538 7398 586622 7634
rect 586858 7398 586890 7634
rect 582294 -1542 582326 -1306
rect 582562 -1542 582646 -1306
rect 582882 -1542 582914 -1306
rect 582294 -1626 582914 -1542
rect 582294 -1862 582326 -1626
rect 582562 -1862 582646 -1626
rect 582882 -1862 582914 -1626
rect 582294 -7654 582914 -1862
rect 586270 -1306 586890 7398
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 696454 587850 706202
rect 587230 696218 587262 696454
rect 587498 696218 587582 696454
rect 587818 696218 587850 696454
rect 587230 696134 587850 696218
rect 587230 695898 587262 696134
rect 587498 695898 587582 696134
rect 587818 695898 587850 696134
rect 587230 660454 587850 695898
rect 587230 660218 587262 660454
rect 587498 660218 587582 660454
rect 587818 660218 587850 660454
rect 587230 660134 587850 660218
rect 587230 659898 587262 660134
rect 587498 659898 587582 660134
rect 587818 659898 587850 660134
rect 587230 624454 587850 659898
rect 587230 624218 587262 624454
rect 587498 624218 587582 624454
rect 587818 624218 587850 624454
rect 587230 624134 587850 624218
rect 587230 623898 587262 624134
rect 587498 623898 587582 624134
rect 587818 623898 587850 624134
rect 587230 588454 587850 623898
rect 587230 588218 587262 588454
rect 587498 588218 587582 588454
rect 587818 588218 587850 588454
rect 587230 588134 587850 588218
rect 587230 587898 587262 588134
rect 587498 587898 587582 588134
rect 587818 587898 587850 588134
rect 587230 552454 587850 587898
rect 587230 552218 587262 552454
rect 587498 552218 587582 552454
rect 587818 552218 587850 552454
rect 587230 552134 587850 552218
rect 587230 551898 587262 552134
rect 587498 551898 587582 552134
rect 587818 551898 587850 552134
rect 587230 516454 587850 551898
rect 587230 516218 587262 516454
rect 587498 516218 587582 516454
rect 587818 516218 587850 516454
rect 587230 516134 587850 516218
rect 587230 515898 587262 516134
rect 587498 515898 587582 516134
rect 587818 515898 587850 516134
rect 587230 480454 587850 515898
rect 587230 480218 587262 480454
rect 587498 480218 587582 480454
rect 587818 480218 587850 480454
rect 587230 480134 587850 480218
rect 587230 479898 587262 480134
rect 587498 479898 587582 480134
rect 587818 479898 587850 480134
rect 587230 444454 587850 479898
rect 587230 444218 587262 444454
rect 587498 444218 587582 444454
rect 587818 444218 587850 444454
rect 587230 444134 587850 444218
rect 587230 443898 587262 444134
rect 587498 443898 587582 444134
rect 587818 443898 587850 444134
rect 587230 408454 587850 443898
rect 587230 408218 587262 408454
rect 587498 408218 587582 408454
rect 587818 408218 587850 408454
rect 587230 408134 587850 408218
rect 587230 407898 587262 408134
rect 587498 407898 587582 408134
rect 587818 407898 587850 408134
rect 587230 372454 587850 407898
rect 587230 372218 587262 372454
rect 587498 372218 587582 372454
rect 587818 372218 587850 372454
rect 587230 372134 587850 372218
rect 587230 371898 587262 372134
rect 587498 371898 587582 372134
rect 587818 371898 587850 372134
rect 587230 336454 587850 371898
rect 587230 336218 587262 336454
rect 587498 336218 587582 336454
rect 587818 336218 587850 336454
rect 587230 336134 587850 336218
rect 587230 335898 587262 336134
rect 587498 335898 587582 336134
rect 587818 335898 587850 336134
rect 587230 300454 587850 335898
rect 587230 300218 587262 300454
rect 587498 300218 587582 300454
rect 587818 300218 587850 300454
rect 587230 300134 587850 300218
rect 587230 299898 587262 300134
rect 587498 299898 587582 300134
rect 587818 299898 587850 300134
rect 587230 264454 587850 299898
rect 587230 264218 587262 264454
rect 587498 264218 587582 264454
rect 587818 264218 587850 264454
rect 587230 264134 587850 264218
rect 587230 263898 587262 264134
rect 587498 263898 587582 264134
rect 587818 263898 587850 264134
rect 587230 228454 587850 263898
rect 587230 228218 587262 228454
rect 587498 228218 587582 228454
rect 587818 228218 587850 228454
rect 587230 228134 587850 228218
rect 587230 227898 587262 228134
rect 587498 227898 587582 228134
rect 587818 227898 587850 228134
rect 587230 192454 587850 227898
rect 587230 192218 587262 192454
rect 587498 192218 587582 192454
rect 587818 192218 587850 192454
rect 587230 192134 587850 192218
rect 587230 191898 587262 192134
rect 587498 191898 587582 192134
rect 587818 191898 587850 192134
rect 587230 156454 587850 191898
rect 587230 156218 587262 156454
rect 587498 156218 587582 156454
rect 587818 156218 587850 156454
rect 587230 156134 587850 156218
rect 587230 155898 587262 156134
rect 587498 155898 587582 156134
rect 587818 155898 587850 156134
rect 587230 120454 587850 155898
rect 587230 120218 587262 120454
rect 587498 120218 587582 120454
rect 587818 120218 587850 120454
rect 587230 120134 587850 120218
rect 587230 119898 587262 120134
rect 587498 119898 587582 120134
rect 587818 119898 587850 120134
rect 587230 84454 587850 119898
rect 587230 84218 587262 84454
rect 587498 84218 587582 84454
rect 587818 84218 587850 84454
rect 587230 84134 587850 84218
rect 587230 83898 587262 84134
rect 587498 83898 587582 84134
rect 587818 83898 587850 84134
rect 587230 48454 587850 83898
rect 587230 48218 587262 48454
rect 587498 48218 587582 48454
rect 587818 48218 587850 48454
rect 587230 48134 587850 48218
rect 587230 47898 587262 48134
rect 587498 47898 587582 48134
rect 587818 47898 587850 48134
rect 587230 12454 587850 47898
rect 587230 12218 587262 12454
rect 587498 12218 587582 12454
rect 587818 12218 587850 12454
rect 587230 12134 587850 12218
rect 587230 11898 587262 12134
rect 587498 11898 587582 12134
rect 587818 11898 587850 12134
rect 587230 -2266 587850 11898
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 700954 588810 707162
rect 588190 700718 588222 700954
rect 588458 700718 588542 700954
rect 588778 700718 588810 700954
rect 588190 700634 588810 700718
rect 588190 700398 588222 700634
rect 588458 700398 588542 700634
rect 588778 700398 588810 700634
rect 588190 664954 588810 700398
rect 588190 664718 588222 664954
rect 588458 664718 588542 664954
rect 588778 664718 588810 664954
rect 588190 664634 588810 664718
rect 588190 664398 588222 664634
rect 588458 664398 588542 664634
rect 588778 664398 588810 664634
rect 588190 628954 588810 664398
rect 588190 628718 588222 628954
rect 588458 628718 588542 628954
rect 588778 628718 588810 628954
rect 588190 628634 588810 628718
rect 588190 628398 588222 628634
rect 588458 628398 588542 628634
rect 588778 628398 588810 628634
rect 588190 592954 588810 628398
rect 588190 592718 588222 592954
rect 588458 592718 588542 592954
rect 588778 592718 588810 592954
rect 588190 592634 588810 592718
rect 588190 592398 588222 592634
rect 588458 592398 588542 592634
rect 588778 592398 588810 592634
rect 588190 556954 588810 592398
rect 588190 556718 588222 556954
rect 588458 556718 588542 556954
rect 588778 556718 588810 556954
rect 588190 556634 588810 556718
rect 588190 556398 588222 556634
rect 588458 556398 588542 556634
rect 588778 556398 588810 556634
rect 588190 520954 588810 556398
rect 588190 520718 588222 520954
rect 588458 520718 588542 520954
rect 588778 520718 588810 520954
rect 588190 520634 588810 520718
rect 588190 520398 588222 520634
rect 588458 520398 588542 520634
rect 588778 520398 588810 520634
rect 588190 484954 588810 520398
rect 588190 484718 588222 484954
rect 588458 484718 588542 484954
rect 588778 484718 588810 484954
rect 588190 484634 588810 484718
rect 588190 484398 588222 484634
rect 588458 484398 588542 484634
rect 588778 484398 588810 484634
rect 588190 448954 588810 484398
rect 588190 448718 588222 448954
rect 588458 448718 588542 448954
rect 588778 448718 588810 448954
rect 588190 448634 588810 448718
rect 588190 448398 588222 448634
rect 588458 448398 588542 448634
rect 588778 448398 588810 448634
rect 588190 412954 588810 448398
rect 588190 412718 588222 412954
rect 588458 412718 588542 412954
rect 588778 412718 588810 412954
rect 588190 412634 588810 412718
rect 588190 412398 588222 412634
rect 588458 412398 588542 412634
rect 588778 412398 588810 412634
rect 588190 376954 588810 412398
rect 588190 376718 588222 376954
rect 588458 376718 588542 376954
rect 588778 376718 588810 376954
rect 588190 376634 588810 376718
rect 588190 376398 588222 376634
rect 588458 376398 588542 376634
rect 588778 376398 588810 376634
rect 588190 340954 588810 376398
rect 588190 340718 588222 340954
rect 588458 340718 588542 340954
rect 588778 340718 588810 340954
rect 588190 340634 588810 340718
rect 588190 340398 588222 340634
rect 588458 340398 588542 340634
rect 588778 340398 588810 340634
rect 588190 304954 588810 340398
rect 588190 304718 588222 304954
rect 588458 304718 588542 304954
rect 588778 304718 588810 304954
rect 588190 304634 588810 304718
rect 588190 304398 588222 304634
rect 588458 304398 588542 304634
rect 588778 304398 588810 304634
rect 588190 268954 588810 304398
rect 588190 268718 588222 268954
rect 588458 268718 588542 268954
rect 588778 268718 588810 268954
rect 588190 268634 588810 268718
rect 588190 268398 588222 268634
rect 588458 268398 588542 268634
rect 588778 268398 588810 268634
rect 588190 232954 588810 268398
rect 588190 232718 588222 232954
rect 588458 232718 588542 232954
rect 588778 232718 588810 232954
rect 588190 232634 588810 232718
rect 588190 232398 588222 232634
rect 588458 232398 588542 232634
rect 588778 232398 588810 232634
rect 588190 196954 588810 232398
rect 588190 196718 588222 196954
rect 588458 196718 588542 196954
rect 588778 196718 588810 196954
rect 588190 196634 588810 196718
rect 588190 196398 588222 196634
rect 588458 196398 588542 196634
rect 588778 196398 588810 196634
rect 588190 160954 588810 196398
rect 588190 160718 588222 160954
rect 588458 160718 588542 160954
rect 588778 160718 588810 160954
rect 588190 160634 588810 160718
rect 588190 160398 588222 160634
rect 588458 160398 588542 160634
rect 588778 160398 588810 160634
rect 588190 124954 588810 160398
rect 588190 124718 588222 124954
rect 588458 124718 588542 124954
rect 588778 124718 588810 124954
rect 588190 124634 588810 124718
rect 588190 124398 588222 124634
rect 588458 124398 588542 124634
rect 588778 124398 588810 124634
rect 588190 88954 588810 124398
rect 588190 88718 588222 88954
rect 588458 88718 588542 88954
rect 588778 88718 588810 88954
rect 588190 88634 588810 88718
rect 588190 88398 588222 88634
rect 588458 88398 588542 88634
rect 588778 88398 588810 88634
rect 588190 52954 588810 88398
rect 588190 52718 588222 52954
rect 588458 52718 588542 52954
rect 588778 52718 588810 52954
rect 588190 52634 588810 52718
rect 588190 52398 588222 52634
rect 588458 52398 588542 52634
rect 588778 52398 588810 52634
rect 588190 16954 588810 52398
rect 588190 16718 588222 16954
rect 588458 16718 588542 16954
rect 588778 16718 588810 16954
rect 588190 16634 588810 16718
rect 588190 16398 588222 16634
rect 588458 16398 588542 16634
rect 588778 16398 588810 16634
rect 588190 -3226 588810 16398
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 669454 589770 708122
rect 589150 669218 589182 669454
rect 589418 669218 589502 669454
rect 589738 669218 589770 669454
rect 589150 669134 589770 669218
rect 589150 668898 589182 669134
rect 589418 668898 589502 669134
rect 589738 668898 589770 669134
rect 589150 633454 589770 668898
rect 589150 633218 589182 633454
rect 589418 633218 589502 633454
rect 589738 633218 589770 633454
rect 589150 633134 589770 633218
rect 589150 632898 589182 633134
rect 589418 632898 589502 633134
rect 589738 632898 589770 633134
rect 589150 597454 589770 632898
rect 589150 597218 589182 597454
rect 589418 597218 589502 597454
rect 589738 597218 589770 597454
rect 589150 597134 589770 597218
rect 589150 596898 589182 597134
rect 589418 596898 589502 597134
rect 589738 596898 589770 597134
rect 589150 561454 589770 596898
rect 589150 561218 589182 561454
rect 589418 561218 589502 561454
rect 589738 561218 589770 561454
rect 589150 561134 589770 561218
rect 589150 560898 589182 561134
rect 589418 560898 589502 561134
rect 589738 560898 589770 561134
rect 589150 525454 589770 560898
rect 589150 525218 589182 525454
rect 589418 525218 589502 525454
rect 589738 525218 589770 525454
rect 589150 525134 589770 525218
rect 589150 524898 589182 525134
rect 589418 524898 589502 525134
rect 589738 524898 589770 525134
rect 589150 489454 589770 524898
rect 589150 489218 589182 489454
rect 589418 489218 589502 489454
rect 589738 489218 589770 489454
rect 589150 489134 589770 489218
rect 589150 488898 589182 489134
rect 589418 488898 589502 489134
rect 589738 488898 589770 489134
rect 589150 453454 589770 488898
rect 589150 453218 589182 453454
rect 589418 453218 589502 453454
rect 589738 453218 589770 453454
rect 589150 453134 589770 453218
rect 589150 452898 589182 453134
rect 589418 452898 589502 453134
rect 589738 452898 589770 453134
rect 589150 417454 589770 452898
rect 589150 417218 589182 417454
rect 589418 417218 589502 417454
rect 589738 417218 589770 417454
rect 589150 417134 589770 417218
rect 589150 416898 589182 417134
rect 589418 416898 589502 417134
rect 589738 416898 589770 417134
rect 589150 381454 589770 416898
rect 589150 381218 589182 381454
rect 589418 381218 589502 381454
rect 589738 381218 589770 381454
rect 589150 381134 589770 381218
rect 589150 380898 589182 381134
rect 589418 380898 589502 381134
rect 589738 380898 589770 381134
rect 589150 345454 589770 380898
rect 589150 345218 589182 345454
rect 589418 345218 589502 345454
rect 589738 345218 589770 345454
rect 589150 345134 589770 345218
rect 589150 344898 589182 345134
rect 589418 344898 589502 345134
rect 589738 344898 589770 345134
rect 589150 309454 589770 344898
rect 589150 309218 589182 309454
rect 589418 309218 589502 309454
rect 589738 309218 589770 309454
rect 589150 309134 589770 309218
rect 589150 308898 589182 309134
rect 589418 308898 589502 309134
rect 589738 308898 589770 309134
rect 589150 273454 589770 308898
rect 589150 273218 589182 273454
rect 589418 273218 589502 273454
rect 589738 273218 589770 273454
rect 589150 273134 589770 273218
rect 589150 272898 589182 273134
rect 589418 272898 589502 273134
rect 589738 272898 589770 273134
rect 589150 237454 589770 272898
rect 589150 237218 589182 237454
rect 589418 237218 589502 237454
rect 589738 237218 589770 237454
rect 589150 237134 589770 237218
rect 589150 236898 589182 237134
rect 589418 236898 589502 237134
rect 589738 236898 589770 237134
rect 589150 201454 589770 236898
rect 589150 201218 589182 201454
rect 589418 201218 589502 201454
rect 589738 201218 589770 201454
rect 589150 201134 589770 201218
rect 589150 200898 589182 201134
rect 589418 200898 589502 201134
rect 589738 200898 589770 201134
rect 589150 165454 589770 200898
rect 589150 165218 589182 165454
rect 589418 165218 589502 165454
rect 589738 165218 589770 165454
rect 589150 165134 589770 165218
rect 589150 164898 589182 165134
rect 589418 164898 589502 165134
rect 589738 164898 589770 165134
rect 589150 129454 589770 164898
rect 589150 129218 589182 129454
rect 589418 129218 589502 129454
rect 589738 129218 589770 129454
rect 589150 129134 589770 129218
rect 589150 128898 589182 129134
rect 589418 128898 589502 129134
rect 589738 128898 589770 129134
rect 589150 93454 589770 128898
rect 589150 93218 589182 93454
rect 589418 93218 589502 93454
rect 589738 93218 589770 93454
rect 589150 93134 589770 93218
rect 589150 92898 589182 93134
rect 589418 92898 589502 93134
rect 589738 92898 589770 93134
rect 589150 57454 589770 92898
rect 589150 57218 589182 57454
rect 589418 57218 589502 57454
rect 589738 57218 589770 57454
rect 589150 57134 589770 57218
rect 589150 56898 589182 57134
rect 589418 56898 589502 57134
rect 589738 56898 589770 57134
rect 589150 21454 589770 56898
rect 589150 21218 589182 21454
rect 589418 21218 589502 21454
rect 589738 21218 589770 21454
rect 589150 21134 589770 21218
rect 589150 20898 589182 21134
rect 589418 20898 589502 21134
rect 589738 20898 589770 21134
rect 589150 -4186 589770 20898
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 673954 590730 709082
rect 590110 673718 590142 673954
rect 590378 673718 590462 673954
rect 590698 673718 590730 673954
rect 590110 673634 590730 673718
rect 590110 673398 590142 673634
rect 590378 673398 590462 673634
rect 590698 673398 590730 673634
rect 590110 637954 590730 673398
rect 590110 637718 590142 637954
rect 590378 637718 590462 637954
rect 590698 637718 590730 637954
rect 590110 637634 590730 637718
rect 590110 637398 590142 637634
rect 590378 637398 590462 637634
rect 590698 637398 590730 637634
rect 590110 601954 590730 637398
rect 590110 601718 590142 601954
rect 590378 601718 590462 601954
rect 590698 601718 590730 601954
rect 590110 601634 590730 601718
rect 590110 601398 590142 601634
rect 590378 601398 590462 601634
rect 590698 601398 590730 601634
rect 590110 565954 590730 601398
rect 590110 565718 590142 565954
rect 590378 565718 590462 565954
rect 590698 565718 590730 565954
rect 590110 565634 590730 565718
rect 590110 565398 590142 565634
rect 590378 565398 590462 565634
rect 590698 565398 590730 565634
rect 590110 529954 590730 565398
rect 590110 529718 590142 529954
rect 590378 529718 590462 529954
rect 590698 529718 590730 529954
rect 590110 529634 590730 529718
rect 590110 529398 590142 529634
rect 590378 529398 590462 529634
rect 590698 529398 590730 529634
rect 590110 493954 590730 529398
rect 590110 493718 590142 493954
rect 590378 493718 590462 493954
rect 590698 493718 590730 493954
rect 590110 493634 590730 493718
rect 590110 493398 590142 493634
rect 590378 493398 590462 493634
rect 590698 493398 590730 493634
rect 590110 457954 590730 493398
rect 590110 457718 590142 457954
rect 590378 457718 590462 457954
rect 590698 457718 590730 457954
rect 590110 457634 590730 457718
rect 590110 457398 590142 457634
rect 590378 457398 590462 457634
rect 590698 457398 590730 457634
rect 590110 421954 590730 457398
rect 590110 421718 590142 421954
rect 590378 421718 590462 421954
rect 590698 421718 590730 421954
rect 590110 421634 590730 421718
rect 590110 421398 590142 421634
rect 590378 421398 590462 421634
rect 590698 421398 590730 421634
rect 590110 385954 590730 421398
rect 590110 385718 590142 385954
rect 590378 385718 590462 385954
rect 590698 385718 590730 385954
rect 590110 385634 590730 385718
rect 590110 385398 590142 385634
rect 590378 385398 590462 385634
rect 590698 385398 590730 385634
rect 590110 349954 590730 385398
rect 590110 349718 590142 349954
rect 590378 349718 590462 349954
rect 590698 349718 590730 349954
rect 590110 349634 590730 349718
rect 590110 349398 590142 349634
rect 590378 349398 590462 349634
rect 590698 349398 590730 349634
rect 590110 313954 590730 349398
rect 590110 313718 590142 313954
rect 590378 313718 590462 313954
rect 590698 313718 590730 313954
rect 590110 313634 590730 313718
rect 590110 313398 590142 313634
rect 590378 313398 590462 313634
rect 590698 313398 590730 313634
rect 590110 277954 590730 313398
rect 590110 277718 590142 277954
rect 590378 277718 590462 277954
rect 590698 277718 590730 277954
rect 590110 277634 590730 277718
rect 590110 277398 590142 277634
rect 590378 277398 590462 277634
rect 590698 277398 590730 277634
rect 590110 241954 590730 277398
rect 590110 241718 590142 241954
rect 590378 241718 590462 241954
rect 590698 241718 590730 241954
rect 590110 241634 590730 241718
rect 590110 241398 590142 241634
rect 590378 241398 590462 241634
rect 590698 241398 590730 241634
rect 590110 205954 590730 241398
rect 590110 205718 590142 205954
rect 590378 205718 590462 205954
rect 590698 205718 590730 205954
rect 590110 205634 590730 205718
rect 590110 205398 590142 205634
rect 590378 205398 590462 205634
rect 590698 205398 590730 205634
rect 590110 169954 590730 205398
rect 590110 169718 590142 169954
rect 590378 169718 590462 169954
rect 590698 169718 590730 169954
rect 590110 169634 590730 169718
rect 590110 169398 590142 169634
rect 590378 169398 590462 169634
rect 590698 169398 590730 169634
rect 590110 133954 590730 169398
rect 590110 133718 590142 133954
rect 590378 133718 590462 133954
rect 590698 133718 590730 133954
rect 590110 133634 590730 133718
rect 590110 133398 590142 133634
rect 590378 133398 590462 133634
rect 590698 133398 590730 133634
rect 590110 97954 590730 133398
rect 590110 97718 590142 97954
rect 590378 97718 590462 97954
rect 590698 97718 590730 97954
rect 590110 97634 590730 97718
rect 590110 97398 590142 97634
rect 590378 97398 590462 97634
rect 590698 97398 590730 97634
rect 590110 61954 590730 97398
rect 590110 61718 590142 61954
rect 590378 61718 590462 61954
rect 590698 61718 590730 61954
rect 590110 61634 590730 61718
rect 590110 61398 590142 61634
rect 590378 61398 590462 61634
rect 590698 61398 590730 61634
rect 590110 25954 590730 61398
rect 590110 25718 590142 25954
rect 590378 25718 590462 25954
rect 590698 25718 590730 25954
rect 590110 25634 590730 25718
rect 590110 25398 590142 25634
rect 590378 25398 590462 25634
rect 590698 25398 590730 25634
rect 590110 -5146 590730 25398
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 678454 591690 710042
rect 591070 678218 591102 678454
rect 591338 678218 591422 678454
rect 591658 678218 591690 678454
rect 591070 678134 591690 678218
rect 591070 677898 591102 678134
rect 591338 677898 591422 678134
rect 591658 677898 591690 678134
rect 591070 642454 591690 677898
rect 591070 642218 591102 642454
rect 591338 642218 591422 642454
rect 591658 642218 591690 642454
rect 591070 642134 591690 642218
rect 591070 641898 591102 642134
rect 591338 641898 591422 642134
rect 591658 641898 591690 642134
rect 591070 606454 591690 641898
rect 591070 606218 591102 606454
rect 591338 606218 591422 606454
rect 591658 606218 591690 606454
rect 591070 606134 591690 606218
rect 591070 605898 591102 606134
rect 591338 605898 591422 606134
rect 591658 605898 591690 606134
rect 591070 570454 591690 605898
rect 591070 570218 591102 570454
rect 591338 570218 591422 570454
rect 591658 570218 591690 570454
rect 591070 570134 591690 570218
rect 591070 569898 591102 570134
rect 591338 569898 591422 570134
rect 591658 569898 591690 570134
rect 591070 534454 591690 569898
rect 591070 534218 591102 534454
rect 591338 534218 591422 534454
rect 591658 534218 591690 534454
rect 591070 534134 591690 534218
rect 591070 533898 591102 534134
rect 591338 533898 591422 534134
rect 591658 533898 591690 534134
rect 591070 498454 591690 533898
rect 591070 498218 591102 498454
rect 591338 498218 591422 498454
rect 591658 498218 591690 498454
rect 591070 498134 591690 498218
rect 591070 497898 591102 498134
rect 591338 497898 591422 498134
rect 591658 497898 591690 498134
rect 591070 462454 591690 497898
rect 591070 462218 591102 462454
rect 591338 462218 591422 462454
rect 591658 462218 591690 462454
rect 591070 462134 591690 462218
rect 591070 461898 591102 462134
rect 591338 461898 591422 462134
rect 591658 461898 591690 462134
rect 591070 426454 591690 461898
rect 591070 426218 591102 426454
rect 591338 426218 591422 426454
rect 591658 426218 591690 426454
rect 591070 426134 591690 426218
rect 591070 425898 591102 426134
rect 591338 425898 591422 426134
rect 591658 425898 591690 426134
rect 591070 390454 591690 425898
rect 591070 390218 591102 390454
rect 591338 390218 591422 390454
rect 591658 390218 591690 390454
rect 591070 390134 591690 390218
rect 591070 389898 591102 390134
rect 591338 389898 591422 390134
rect 591658 389898 591690 390134
rect 591070 354454 591690 389898
rect 591070 354218 591102 354454
rect 591338 354218 591422 354454
rect 591658 354218 591690 354454
rect 591070 354134 591690 354218
rect 591070 353898 591102 354134
rect 591338 353898 591422 354134
rect 591658 353898 591690 354134
rect 591070 318454 591690 353898
rect 591070 318218 591102 318454
rect 591338 318218 591422 318454
rect 591658 318218 591690 318454
rect 591070 318134 591690 318218
rect 591070 317898 591102 318134
rect 591338 317898 591422 318134
rect 591658 317898 591690 318134
rect 591070 282454 591690 317898
rect 591070 282218 591102 282454
rect 591338 282218 591422 282454
rect 591658 282218 591690 282454
rect 591070 282134 591690 282218
rect 591070 281898 591102 282134
rect 591338 281898 591422 282134
rect 591658 281898 591690 282134
rect 591070 246454 591690 281898
rect 591070 246218 591102 246454
rect 591338 246218 591422 246454
rect 591658 246218 591690 246454
rect 591070 246134 591690 246218
rect 591070 245898 591102 246134
rect 591338 245898 591422 246134
rect 591658 245898 591690 246134
rect 591070 210454 591690 245898
rect 591070 210218 591102 210454
rect 591338 210218 591422 210454
rect 591658 210218 591690 210454
rect 591070 210134 591690 210218
rect 591070 209898 591102 210134
rect 591338 209898 591422 210134
rect 591658 209898 591690 210134
rect 591070 174454 591690 209898
rect 591070 174218 591102 174454
rect 591338 174218 591422 174454
rect 591658 174218 591690 174454
rect 591070 174134 591690 174218
rect 591070 173898 591102 174134
rect 591338 173898 591422 174134
rect 591658 173898 591690 174134
rect 591070 138454 591690 173898
rect 591070 138218 591102 138454
rect 591338 138218 591422 138454
rect 591658 138218 591690 138454
rect 591070 138134 591690 138218
rect 591070 137898 591102 138134
rect 591338 137898 591422 138134
rect 591658 137898 591690 138134
rect 591070 102454 591690 137898
rect 591070 102218 591102 102454
rect 591338 102218 591422 102454
rect 591658 102218 591690 102454
rect 591070 102134 591690 102218
rect 591070 101898 591102 102134
rect 591338 101898 591422 102134
rect 591658 101898 591690 102134
rect 591070 66454 591690 101898
rect 591070 66218 591102 66454
rect 591338 66218 591422 66454
rect 591658 66218 591690 66454
rect 591070 66134 591690 66218
rect 591070 65898 591102 66134
rect 591338 65898 591422 66134
rect 591658 65898 591690 66134
rect 591070 30454 591690 65898
rect 591070 30218 591102 30454
rect 591338 30218 591422 30454
rect 591658 30218 591690 30454
rect 591070 30134 591690 30218
rect 591070 29898 591102 30134
rect 591338 29898 591422 30134
rect 591658 29898 591690 30134
rect 591070 -6106 591690 29898
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 682954 592650 711002
rect 592030 682718 592062 682954
rect 592298 682718 592382 682954
rect 592618 682718 592650 682954
rect 592030 682634 592650 682718
rect 592030 682398 592062 682634
rect 592298 682398 592382 682634
rect 592618 682398 592650 682634
rect 592030 646954 592650 682398
rect 592030 646718 592062 646954
rect 592298 646718 592382 646954
rect 592618 646718 592650 646954
rect 592030 646634 592650 646718
rect 592030 646398 592062 646634
rect 592298 646398 592382 646634
rect 592618 646398 592650 646634
rect 592030 610954 592650 646398
rect 592030 610718 592062 610954
rect 592298 610718 592382 610954
rect 592618 610718 592650 610954
rect 592030 610634 592650 610718
rect 592030 610398 592062 610634
rect 592298 610398 592382 610634
rect 592618 610398 592650 610634
rect 592030 574954 592650 610398
rect 592030 574718 592062 574954
rect 592298 574718 592382 574954
rect 592618 574718 592650 574954
rect 592030 574634 592650 574718
rect 592030 574398 592062 574634
rect 592298 574398 592382 574634
rect 592618 574398 592650 574634
rect 592030 538954 592650 574398
rect 592030 538718 592062 538954
rect 592298 538718 592382 538954
rect 592618 538718 592650 538954
rect 592030 538634 592650 538718
rect 592030 538398 592062 538634
rect 592298 538398 592382 538634
rect 592618 538398 592650 538634
rect 592030 502954 592650 538398
rect 592030 502718 592062 502954
rect 592298 502718 592382 502954
rect 592618 502718 592650 502954
rect 592030 502634 592650 502718
rect 592030 502398 592062 502634
rect 592298 502398 592382 502634
rect 592618 502398 592650 502634
rect 592030 466954 592650 502398
rect 592030 466718 592062 466954
rect 592298 466718 592382 466954
rect 592618 466718 592650 466954
rect 592030 466634 592650 466718
rect 592030 466398 592062 466634
rect 592298 466398 592382 466634
rect 592618 466398 592650 466634
rect 592030 430954 592650 466398
rect 592030 430718 592062 430954
rect 592298 430718 592382 430954
rect 592618 430718 592650 430954
rect 592030 430634 592650 430718
rect 592030 430398 592062 430634
rect 592298 430398 592382 430634
rect 592618 430398 592650 430634
rect 592030 394954 592650 430398
rect 592030 394718 592062 394954
rect 592298 394718 592382 394954
rect 592618 394718 592650 394954
rect 592030 394634 592650 394718
rect 592030 394398 592062 394634
rect 592298 394398 592382 394634
rect 592618 394398 592650 394634
rect 592030 358954 592650 394398
rect 592030 358718 592062 358954
rect 592298 358718 592382 358954
rect 592618 358718 592650 358954
rect 592030 358634 592650 358718
rect 592030 358398 592062 358634
rect 592298 358398 592382 358634
rect 592618 358398 592650 358634
rect 592030 322954 592650 358398
rect 592030 322718 592062 322954
rect 592298 322718 592382 322954
rect 592618 322718 592650 322954
rect 592030 322634 592650 322718
rect 592030 322398 592062 322634
rect 592298 322398 592382 322634
rect 592618 322398 592650 322634
rect 592030 286954 592650 322398
rect 592030 286718 592062 286954
rect 592298 286718 592382 286954
rect 592618 286718 592650 286954
rect 592030 286634 592650 286718
rect 592030 286398 592062 286634
rect 592298 286398 592382 286634
rect 592618 286398 592650 286634
rect 592030 250954 592650 286398
rect 592030 250718 592062 250954
rect 592298 250718 592382 250954
rect 592618 250718 592650 250954
rect 592030 250634 592650 250718
rect 592030 250398 592062 250634
rect 592298 250398 592382 250634
rect 592618 250398 592650 250634
rect 592030 214954 592650 250398
rect 592030 214718 592062 214954
rect 592298 214718 592382 214954
rect 592618 214718 592650 214954
rect 592030 214634 592650 214718
rect 592030 214398 592062 214634
rect 592298 214398 592382 214634
rect 592618 214398 592650 214634
rect 592030 178954 592650 214398
rect 592030 178718 592062 178954
rect 592298 178718 592382 178954
rect 592618 178718 592650 178954
rect 592030 178634 592650 178718
rect 592030 178398 592062 178634
rect 592298 178398 592382 178634
rect 592618 178398 592650 178634
rect 592030 142954 592650 178398
rect 592030 142718 592062 142954
rect 592298 142718 592382 142954
rect 592618 142718 592650 142954
rect 592030 142634 592650 142718
rect 592030 142398 592062 142634
rect 592298 142398 592382 142634
rect 592618 142398 592650 142634
rect 592030 106954 592650 142398
rect 592030 106718 592062 106954
rect 592298 106718 592382 106954
rect 592618 106718 592650 106954
rect 592030 106634 592650 106718
rect 592030 106398 592062 106634
rect 592298 106398 592382 106634
rect 592618 106398 592650 106634
rect 592030 70954 592650 106398
rect 592030 70718 592062 70954
rect 592298 70718 592382 70954
rect 592618 70718 592650 70954
rect 592030 70634 592650 70718
rect 592030 70398 592062 70634
rect 592298 70398 592382 70634
rect 592618 70398 592650 70634
rect 592030 34954 592650 70398
rect 592030 34718 592062 34954
rect 592298 34718 592382 34954
rect 592618 34718 592650 34954
rect 592030 34634 592650 34718
rect 592030 34398 592062 34634
rect 592298 34398 592382 34634
rect 592618 34398 592650 34634
rect 592030 -7066 592650 34398
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 682718 -8458 682954
rect -8374 682718 -8138 682954
rect -8694 682398 -8458 682634
rect -8374 682398 -8138 682634
rect -8694 646718 -8458 646954
rect -8374 646718 -8138 646954
rect -8694 646398 -8458 646634
rect -8374 646398 -8138 646634
rect -8694 610718 -8458 610954
rect -8374 610718 -8138 610954
rect -8694 610398 -8458 610634
rect -8374 610398 -8138 610634
rect -8694 574718 -8458 574954
rect -8374 574718 -8138 574954
rect -8694 574398 -8458 574634
rect -8374 574398 -8138 574634
rect -8694 538718 -8458 538954
rect -8374 538718 -8138 538954
rect -8694 538398 -8458 538634
rect -8374 538398 -8138 538634
rect -8694 502718 -8458 502954
rect -8374 502718 -8138 502954
rect -8694 502398 -8458 502634
rect -8374 502398 -8138 502634
rect -8694 466718 -8458 466954
rect -8374 466718 -8138 466954
rect -8694 466398 -8458 466634
rect -8374 466398 -8138 466634
rect -8694 430718 -8458 430954
rect -8374 430718 -8138 430954
rect -8694 430398 -8458 430634
rect -8374 430398 -8138 430634
rect -8694 394718 -8458 394954
rect -8374 394718 -8138 394954
rect -8694 394398 -8458 394634
rect -8374 394398 -8138 394634
rect -8694 358718 -8458 358954
rect -8374 358718 -8138 358954
rect -8694 358398 -8458 358634
rect -8374 358398 -8138 358634
rect -8694 322718 -8458 322954
rect -8374 322718 -8138 322954
rect -8694 322398 -8458 322634
rect -8374 322398 -8138 322634
rect -8694 286718 -8458 286954
rect -8374 286718 -8138 286954
rect -8694 286398 -8458 286634
rect -8374 286398 -8138 286634
rect -8694 250718 -8458 250954
rect -8374 250718 -8138 250954
rect -8694 250398 -8458 250634
rect -8374 250398 -8138 250634
rect -8694 214718 -8458 214954
rect -8374 214718 -8138 214954
rect -8694 214398 -8458 214634
rect -8374 214398 -8138 214634
rect -8694 178718 -8458 178954
rect -8374 178718 -8138 178954
rect -8694 178398 -8458 178634
rect -8374 178398 -8138 178634
rect -8694 142718 -8458 142954
rect -8374 142718 -8138 142954
rect -8694 142398 -8458 142634
rect -8374 142398 -8138 142634
rect -8694 106718 -8458 106954
rect -8374 106718 -8138 106954
rect -8694 106398 -8458 106634
rect -8374 106398 -8138 106634
rect -8694 70718 -8458 70954
rect -8374 70718 -8138 70954
rect -8694 70398 -8458 70634
rect -8374 70398 -8138 70634
rect -8694 34718 -8458 34954
rect -8374 34718 -8138 34954
rect -8694 34398 -8458 34634
rect -8374 34398 -8138 34634
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect -7734 678218 -7498 678454
rect -7414 678218 -7178 678454
rect -7734 677898 -7498 678134
rect -7414 677898 -7178 678134
rect -7734 642218 -7498 642454
rect -7414 642218 -7178 642454
rect -7734 641898 -7498 642134
rect -7414 641898 -7178 642134
rect -7734 606218 -7498 606454
rect -7414 606218 -7178 606454
rect -7734 605898 -7498 606134
rect -7414 605898 -7178 606134
rect -7734 570218 -7498 570454
rect -7414 570218 -7178 570454
rect -7734 569898 -7498 570134
rect -7414 569898 -7178 570134
rect -7734 534218 -7498 534454
rect -7414 534218 -7178 534454
rect -7734 533898 -7498 534134
rect -7414 533898 -7178 534134
rect -7734 498218 -7498 498454
rect -7414 498218 -7178 498454
rect -7734 497898 -7498 498134
rect -7414 497898 -7178 498134
rect -7734 462218 -7498 462454
rect -7414 462218 -7178 462454
rect -7734 461898 -7498 462134
rect -7414 461898 -7178 462134
rect -7734 426218 -7498 426454
rect -7414 426218 -7178 426454
rect -7734 425898 -7498 426134
rect -7414 425898 -7178 426134
rect -7734 390218 -7498 390454
rect -7414 390218 -7178 390454
rect -7734 389898 -7498 390134
rect -7414 389898 -7178 390134
rect -7734 354218 -7498 354454
rect -7414 354218 -7178 354454
rect -7734 353898 -7498 354134
rect -7414 353898 -7178 354134
rect -7734 318218 -7498 318454
rect -7414 318218 -7178 318454
rect -7734 317898 -7498 318134
rect -7414 317898 -7178 318134
rect -7734 282218 -7498 282454
rect -7414 282218 -7178 282454
rect -7734 281898 -7498 282134
rect -7414 281898 -7178 282134
rect -7734 246218 -7498 246454
rect -7414 246218 -7178 246454
rect -7734 245898 -7498 246134
rect -7414 245898 -7178 246134
rect -7734 210218 -7498 210454
rect -7414 210218 -7178 210454
rect -7734 209898 -7498 210134
rect -7414 209898 -7178 210134
rect -7734 174218 -7498 174454
rect -7414 174218 -7178 174454
rect -7734 173898 -7498 174134
rect -7414 173898 -7178 174134
rect -7734 138218 -7498 138454
rect -7414 138218 -7178 138454
rect -7734 137898 -7498 138134
rect -7414 137898 -7178 138134
rect -7734 102218 -7498 102454
rect -7414 102218 -7178 102454
rect -7734 101898 -7498 102134
rect -7414 101898 -7178 102134
rect -7734 66218 -7498 66454
rect -7414 66218 -7178 66454
rect -7734 65898 -7498 66134
rect -7414 65898 -7178 66134
rect -7734 30218 -7498 30454
rect -7414 30218 -7178 30454
rect -7734 29898 -7498 30134
rect -7414 29898 -7178 30134
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 673718 -6538 673954
rect -6454 673718 -6218 673954
rect -6774 673398 -6538 673634
rect -6454 673398 -6218 673634
rect -6774 637718 -6538 637954
rect -6454 637718 -6218 637954
rect -6774 637398 -6538 637634
rect -6454 637398 -6218 637634
rect -6774 601718 -6538 601954
rect -6454 601718 -6218 601954
rect -6774 601398 -6538 601634
rect -6454 601398 -6218 601634
rect -6774 565718 -6538 565954
rect -6454 565718 -6218 565954
rect -6774 565398 -6538 565634
rect -6454 565398 -6218 565634
rect -6774 529718 -6538 529954
rect -6454 529718 -6218 529954
rect -6774 529398 -6538 529634
rect -6454 529398 -6218 529634
rect -6774 493718 -6538 493954
rect -6454 493718 -6218 493954
rect -6774 493398 -6538 493634
rect -6454 493398 -6218 493634
rect -6774 457718 -6538 457954
rect -6454 457718 -6218 457954
rect -6774 457398 -6538 457634
rect -6454 457398 -6218 457634
rect -6774 421718 -6538 421954
rect -6454 421718 -6218 421954
rect -6774 421398 -6538 421634
rect -6454 421398 -6218 421634
rect -6774 385718 -6538 385954
rect -6454 385718 -6218 385954
rect -6774 385398 -6538 385634
rect -6454 385398 -6218 385634
rect -6774 349718 -6538 349954
rect -6454 349718 -6218 349954
rect -6774 349398 -6538 349634
rect -6454 349398 -6218 349634
rect -6774 313718 -6538 313954
rect -6454 313718 -6218 313954
rect -6774 313398 -6538 313634
rect -6454 313398 -6218 313634
rect -6774 277718 -6538 277954
rect -6454 277718 -6218 277954
rect -6774 277398 -6538 277634
rect -6454 277398 -6218 277634
rect -6774 241718 -6538 241954
rect -6454 241718 -6218 241954
rect -6774 241398 -6538 241634
rect -6454 241398 -6218 241634
rect -6774 205718 -6538 205954
rect -6454 205718 -6218 205954
rect -6774 205398 -6538 205634
rect -6454 205398 -6218 205634
rect -6774 169718 -6538 169954
rect -6454 169718 -6218 169954
rect -6774 169398 -6538 169634
rect -6454 169398 -6218 169634
rect -6774 133718 -6538 133954
rect -6454 133718 -6218 133954
rect -6774 133398 -6538 133634
rect -6454 133398 -6218 133634
rect -6774 97718 -6538 97954
rect -6454 97718 -6218 97954
rect -6774 97398 -6538 97634
rect -6454 97398 -6218 97634
rect -6774 61718 -6538 61954
rect -6454 61718 -6218 61954
rect -6774 61398 -6538 61634
rect -6454 61398 -6218 61634
rect -6774 25718 -6538 25954
rect -6454 25718 -6218 25954
rect -6774 25398 -6538 25634
rect -6454 25398 -6218 25634
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect -5814 669218 -5578 669454
rect -5494 669218 -5258 669454
rect -5814 668898 -5578 669134
rect -5494 668898 -5258 669134
rect -5814 633218 -5578 633454
rect -5494 633218 -5258 633454
rect -5814 632898 -5578 633134
rect -5494 632898 -5258 633134
rect -5814 597218 -5578 597454
rect -5494 597218 -5258 597454
rect -5814 596898 -5578 597134
rect -5494 596898 -5258 597134
rect -5814 561218 -5578 561454
rect -5494 561218 -5258 561454
rect -5814 560898 -5578 561134
rect -5494 560898 -5258 561134
rect -5814 525218 -5578 525454
rect -5494 525218 -5258 525454
rect -5814 524898 -5578 525134
rect -5494 524898 -5258 525134
rect -5814 489218 -5578 489454
rect -5494 489218 -5258 489454
rect -5814 488898 -5578 489134
rect -5494 488898 -5258 489134
rect -5814 453218 -5578 453454
rect -5494 453218 -5258 453454
rect -5814 452898 -5578 453134
rect -5494 452898 -5258 453134
rect -5814 417218 -5578 417454
rect -5494 417218 -5258 417454
rect -5814 416898 -5578 417134
rect -5494 416898 -5258 417134
rect -5814 381218 -5578 381454
rect -5494 381218 -5258 381454
rect -5814 380898 -5578 381134
rect -5494 380898 -5258 381134
rect -5814 345218 -5578 345454
rect -5494 345218 -5258 345454
rect -5814 344898 -5578 345134
rect -5494 344898 -5258 345134
rect -5814 309218 -5578 309454
rect -5494 309218 -5258 309454
rect -5814 308898 -5578 309134
rect -5494 308898 -5258 309134
rect -5814 273218 -5578 273454
rect -5494 273218 -5258 273454
rect -5814 272898 -5578 273134
rect -5494 272898 -5258 273134
rect -5814 237218 -5578 237454
rect -5494 237218 -5258 237454
rect -5814 236898 -5578 237134
rect -5494 236898 -5258 237134
rect -5814 201218 -5578 201454
rect -5494 201218 -5258 201454
rect -5814 200898 -5578 201134
rect -5494 200898 -5258 201134
rect -5814 165218 -5578 165454
rect -5494 165218 -5258 165454
rect -5814 164898 -5578 165134
rect -5494 164898 -5258 165134
rect -5814 129218 -5578 129454
rect -5494 129218 -5258 129454
rect -5814 128898 -5578 129134
rect -5494 128898 -5258 129134
rect -5814 93218 -5578 93454
rect -5494 93218 -5258 93454
rect -5814 92898 -5578 93134
rect -5494 92898 -5258 93134
rect -5814 57218 -5578 57454
rect -5494 57218 -5258 57454
rect -5814 56898 -5578 57134
rect -5494 56898 -5258 57134
rect -5814 21218 -5578 21454
rect -5494 21218 -5258 21454
rect -5814 20898 -5578 21134
rect -5494 20898 -5258 21134
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 700718 -4618 700954
rect -4534 700718 -4298 700954
rect -4854 700398 -4618 700634
rect -4534 700398 -4298 700634
rect -4854 664718 -4618 664954
rect -4534 664718 -4298 664954
rect -4854 664398 -4618 664634
rect -4534 664398 -4298 664634
rect -4854 628718 -4618 628954
rect -4534 628718 -4298 628954
rect -4854 628398 -4618 628634
rect -4534 628398 -4298 628634
rect -4854 592718 -4618 592954
rect -4534 592718 -4298 592954
rect -4854 592398 -4618 592634
rect -4534 592398 -4298 592634
rect -4854 556718 -4618 556954
rect -4534 556718 -4298 556954
rect -4854 556398 -4618 556634
rect -4534 556398 -4298 556634
rect -4854 520718 -4618 520954
rect -4534 520718 -4298 520954
rect -4854 520398 -4618 520634
rect -4534 520398 -4298 520634
rect -4854 484718 -4618 484954
rect -4534 484718 -4298 484954
rect -4854 484398 -4618 484634
rect -4534 484398 -4298 484634
rect -4854 448718 -4618 448954
rect -4534 448718 -4298 448954
rect -4854 448398 -4618 448634
rect -4534 448398 -4298 448634
rect -4854 412718 -4618 412954
rect -4534 412718 -4298 412954
rect -4854 412398 -4618 412634
rect -4534 412398 -4298 412634
rect -4854 376718 -4618 376954
rect -4534 376718 -4298 376954
rect -4854 376398 -4618 376634
rect -4534 376398 -4298 376634
rect -4854 340718 -4618 340954
rect -4534 340718 -4298 340954
rect -4854 340398 -4618 340634
rect -4534 340398 -4298 340634
rect -4854 304718 -4618 304954
rect -4534 304718 -4298 304954
rect -4854 304398 -4618 304634
rect -4534 304398 -4298 304634
rect -4854 268718 -4618 268954
rect -4534 268718 -4298 268954
rect -4854 268398 -4618 268634
rect -4534 268398 -4298 268634
rect -4854 232718 -4618 232954
rect -4534 232718 -4298 232954
rect -4854 232398 -4618 232634
rect -4534 232398 -4298 232634
rect -4854 196718 -4618 196954
rect -4534 196718 -4298 196954
rect -4854 196398 -4618 196634
rect -4534 196398 -4298 196634
rect -4854 160718 -4618 160954
rect -4534 160718 -4298 160954
rect -4854 160398 -4618 160634
rect -4534 160398 -4298 160634
rect -4854 124718 -4618 124954
rect -4534 124718 -4298 124954
rect -4854 124398 -4618 124634
rect -4534 124398 -4298 124634
rect -4854 88718 -4618 88954
rect -4534 88718 -4298 88954
rect -4854 88398 -4618 88634
rect -4534 88398 -4298 88634
rect -4854 52718 -4618 52954
rect -4534 52718 -4298 52954
rect -4854 52398 -4618 52634
rect -4534 52398 -4298 52634
rect -4854 16718 -4618 16954
rect -4534 16718 -4298 16954
rect -4854 16398 -4618 16634
rect -4534 16398 -4298 16634
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect -3894 696218 -3658 696454
rect -3574 696218 -3338 696454
rect -3894 695898 -3658 696134
rect -3574 695898 -3338 696134
rect -3894 660218 -3658 660454
rect -3574 660218 -3338 660454
rect -3894 659898 -3658 660134
rect -3574 659898 -3338 660134
rect -3894 624218 -3658 624454
rect -3574 624218 -3338 624454
rect -3894 623898 -3658 624134
rect -3574 623898 -3338 624134
rect -3894 588218 -3658 588454
rect -3574 588218 -3338 588454
rect -3894 587898 -3658 588134
rect -3574 587898 -3338 588134
rect -3894 552218 -3658 552454
rect -3574 552218 -3338 552454
rect -3894 551898 -3658 552134
rect -3574 551898 -3338 552134
rect -3894 516218 -3658 516454
rect -3574 516218 -3338 516454
rect -3894 515898 -3658 516134
rect -3574 515898 -3338 516134
rect -3894 480218 -3658 480454
rect -3574 480218 -3338 480454
rect -3894 479898 -3658 480134
rect -3574 479898 -3338 480134
rect -3894 444218 -3658 444454
rect -3574 444218 -3338 444454
rect -3894 443898 -3658 444134
rect -3574 443898 -3338 444134
rect -3894 408218 -3658 408454
rect -3574 408218 -3338 408454
rect -3894 407898 -3658 408134
rect -3574 407898 -3338 408134
rect -3894 372218 -3658 372454
rect -3574 372218 -3338 372454
rect -3894 371898 -3658 372134
rect -3574 371898 -3338 372134
rect -3894 336218 -3658 336454
rect -3574 336218 -3338 336454
rect -3894 335898 -3658 336134
rect -3574 335898 -3338 336134
rect -3894 300218 -3658 300454
rect -3574 300218 -3338 300454
rect -3894 299898 -3658 300134
rect -3574 299898 -3338 300134
rect -3894 264218 -3658 264454
rect -3574 264218 -3338 264454
rect -3894 263898 -3658 264134
rect -3574 263898 -3338 264134
rect -3894 228218 -3658 228454
rect -3574 228218 -3338 228454
rect -3894 227898 -3658 228134
rect -3574 227898 -3338 228134
rect -3894 192218 -3658 192454
rect -3574 192218 -3338 192454
rect -3894 191898 -3658 192134
rect -3574 191898 -3338 192134
rect -3894 156218 -3658 156454
rect -3574 156218 -3338 156454
rect -3894 155898 -3658 156134
rect -3574 155898 -3338 156134
rect -3894 120218 -3658 120454
rect -3574 120218 -3338 120454
rect -3894 119898 -3658 120134
rect -3574 119898 -3338 120134
rect -3894 84218 -3658 84454
rect -3574 84218 -3338 84454
rect -3894 83898 -3658 84134
rect -3574 83898 -3338 84134
rect -3894 48218 -3658 48454
rect -3574 48218 -3338 48454
rect -3894 47898 -3658 48134
rect -3574 47898 -3338 48134
rect -3894 12218 -3658 12454
rect -3574 12218 -3338 12454
rect -3894 11898 -3658 12134
rect -3574 11898 -3338 12134
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 691718 -2698 691954
rect -2614 691718 -2378 691954
rect -2934 691398 -2698 691634
rect -2614 691398 -2378 691634
rect -2934 655718 -2698 655954
rect -2614 655718 -2378 655954
rect -2934 655398 -2698 655634
rect -2614 655398 -2378 655634
rect -2934 619718 -2698 619954
rect -2614 619718 -2378 619954
rect -2934 619398 -2698 619634
rect -2614 619398 -2378 619634
rect -2934 583718 -2698 583954
rect -2614 583718 -2378 583954
rect -2934 583398 -2698 583634
rect -2614 583398 -2378 583634
rect -2934 547718 -2698 547954
rect -2614 547718 -2378 547954
rect -2934 547398 -2698 547634
rect -2614 547398 -2378 547634
rect -2934 511718 -2698 511954
rect -2614 511718 -2378 511954
rect -2934 511398 -2698 511634
rect -2614 511398 -2378 511634
rect -2934 475718 -2698 475954
rect -2614 475718 -2378 475954
rect -2934 475398 -2698 475634
rect -2614 475398 -2378 475634
rect -2934 439718 -2698 439954
rect -2614 439718 -2378 439954
rect -2934 439398 -2698 439634
rect -2614 439398 -2378 439634
rect -2934 403718 -2698 403954
rect -2614 403718 -2378 403954
rect -2934 403398 -2698 403634
rect -2614 403398 -2378 403634
rect -2934 367718 -2698 367954
rect -2614 367718 -2378 367954
rect -2934 367398 -2698 367634
rect -2614 367398 -2378 367634
rect -2934 331718 -2698 331954
rect -2614 331718 -2378 331954
rect -2934 331398 -2698 331634
rect -2614 331398 -2378 331634
rect -2934 295718 -2698 295954
rect -2614 295718 -2378 295954
rect -2934 295398 -2698 295634
rect -2614 295398 -2378 295634
rect -2934 259718 -2698 259954
rect -2614 259718 -2378 259954
rect -2934 259398 -2698 259634
rect -2614 259398 -2378 259634
rect -2934 223718 -2698 223954
rect -2614 223718 -2378 223954
rect -2934 223398 -2698 223634
rect -2614 223398 -2378 223634
rect -2934 187718 -2698 187954
rect -2614 187718 -2378 187954
rect -2934 187398 -2698 187634
rect -2614 187398 -2378 187634
rect -2934 151718 -2698 151954
rect -2614 151718 -2378 151954
rect -2934 151398 -2698 151634
rect -2614 151398 -2378 151634
rect -2934 115718 -2698 115954
rect -2614 115718 -2378 115954
rect -2934 115398 -2698 115634
rect -2614 115398 -2378 115634
rect -2934 79718 -2698 79954
rect -2614 79718 -2378 79954
rect -2934 79398 -2698 79634
rect -2614 79398 -2378 79634
rect -2934 43718 -2698 43954
rect -2614 43718 -2378 43954
rect -2934 43398 -2698 43634
rect -2614 43398 -2378 43634
rect -2934 7718 -2698 7954
rect -2614 7718 -2378 7954
rect -2934 7398 -2698 7634
rect -2614 7398 -2378 7634
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 6326 705562 6562 705798
rect 6646 705562 6882 705798
rect 6326 705242 6562 705478
rect 6646 705242 6882 705478
rect 6326 691718 6562 691954
rect 6646 691718 6882 691954
rect 6326 691398 6562 691634
rect 6646 691398 6882 691634
rect 6326 655718 6562 655954
rect 6646 655718 6882 655954
rect 6326 655398 6562 655634
rect 6646 655398 6882 655634
rect 6326 619718 6562 619954
rect 6646 619718 6882 619954
rect 6326 619398 6562 619634
rect 6646 619398 6882 619634
rect 6326 583718 6562 583954
rect 6646 583718 6882 583954
rect 6326 583398 6562 583634
rect 6646 583398 6882 583634
rect 6326 547718 6562 547954
rect 6646 547718 6882 547954
rect 6326 547398 6562 547634
rect 6646 547398 6882 547634
rect 6326 511718 6562 511954
rect 6646 511718 6882 511954
rect 6326 511398 6562 511634
rect 6646 511398 6882 511634
rect 6326 475718 6562 475954
rect 6646 475718 6882 475954
rect 6326 475398 6562 475634
rect 6646 475398 6882 475634
rect 6326 439718 6562 439954
rect 6646 439718 6882 439954
rect 6326 439398 6562 439634
rect 6646 439398 6882 439634
rect 6326 403718 6562 403954
rect 6646 403718 6882 403954
rect 6326 403398 6562 403634
rect 6646 403398 6882 403634
rect 6326 367718 6562 367954
rect 6646 367718 6882 367954
rect 6326 367398 6562 367634
rect 6646 367398 6882 367634
rect 6326 331718 6562 331954
rect 6646 331718 6882 331954
rect 6326 331398 6562 331634
rect 6646 331398 6882 331634
rect 6326 295718 6562 295954
rect 6646 295718 6882 295954
rect 6326 295398 6562 295634
rect 6646 295398 6882 295634
rect 6326 259718 6562 259954
rect 6646 259718 6882 259954
rect 6326 259398 6562 259634
rect 6646 259398 6882 259634
rect 6326 223718 6562 223954
rect 6646 223718 6882 223954
rect 6326 223398 6562 223634
rect 6646 223398 6882 223634
rect 6326 187718 6562 187954
rect 6646 187718 6882 187954
rect 6326 187398 6562 187634
rect 6646 187398 6882 187634
rect 6326 151718 6562 151954
rect 6646 151718 6882 151954
rect 6326 151398 6562 151634
rect 6646 151398 6882 151634
rect 6326 115718 6562 115954
rect 6646 115718 6882 115954
rect 6326 115398 6562 115634
rect 6646 115398 6882 115634
rect 6326 79718 6562 79954
rect 6646 79718 6882 79954
rect 6326 79398 6562 79634
rect 6646 79398 6882 79634
rect 6326 43718 6562 43954
rect 6646 43718 6882 43954
rect 6326 43398 6562 43634
rect 6646 43398 6882 43634
rect 6326 7718 6562 7954
rect 6646 7718 6882 7954
rect 6326 7398 6562 7634
rect 6646 7398 6882 7634
rect 6326 -1542 6562 -1306
rect 6646 -1542 6882 -1306
rect 6326 -1862 6562 -1626
rect 6646 -1862 6882 -1626
rect 10826 706522 11062 706758
rect 11146 706522 11382 706758
rect 10826 706202 11062 706438
rect 11146 706202 11382 706438
rect 10826 696218 11062 696454
rect 11146 696218 11382 696454
rect 10826 695898 11062 696134
rect 11146 695898 11382 696134
rect 10826 660218 11062 660454
rect 11146 660218 11382 660454
rect 10826 659898 11062 660134
rect 11146 659898 11382 660134
rect 10826 624218 11062 624454
rect 11146 624218 11382 624454
rect 10826 623898 11062 624134
rect 11146 623898 11382 624134
rect 10826 588218 11062 588454
rect 11146 588218 11382 588454
rect 10826 587898 11062 588134
rect 11146 587898 11382 588134
rect 10826 552218 11062 552454
rect 11146 552218 11382 552454
rect 10826 551898 11062 552134
rect 11146 551898 11382 552134
rect 10826 516218 11062 516454
rect 11146 516218 11382 516454
rect 10826 515898 11062 516134
rect 11146 515898 11382 516134
rect 10826 480218 11062 480454
rect 11146 480218 11382 480454
rect 10826 479898 11062 480134
rect 11146 479898 11382 480134
rect 10826 444218 11062 444454
rect 11146 444218 11382 444454
rect 10826 443898 11062 444134
rect 11146 443898 11382 444134
rect 10826 408218 11062 408454
rect 11146 408218 11382 408454
rect 10826 407898 11062 408134
rect 11146 407898 11382 408134
rect 10826 372218 11062 372454
rect 11146 372218 11382 372454
rect 10826 371898 11062 372134
rect 11146 371898 11382 372134
rect 10826 336218 11062 336454
rect 11146 336218 11382 336454
rect 10826 335898 11062 336134
rect 11146 335898 11382 336134
rect 10826 300218 11062 300454
rect 11146 300218 11382 300454
rect 10826 299898 11062 300134
rect 11146 299898 11382 300134
rect 10826 264218 11062 264454
rect 11146 264218 11382 264454
rect 10826 263898 11062 264134
rect 11146 263898 11382 264134
rect 10826 228218 11062 228454
rect 11146 228218 11382 228454
rect 10826 227898 11062 228134
rect 11146 227898 11382 228134
rect 10826 192218 11062 192454
rect 11146 192218 11382 192454
rect 10826 191898 11062 192134
rect 11146 191898 11382 192134
rect 10826 156218 11062 156454
rect 11146 156218 11382 156454
rect 10826 155898 11062 156134
rect 11146 155898 11382 156134
rect 10826 120218 11062 120454
rect 11146 120218 11382 120454
rect 10826 119898 11062 120134
rect 11146 119898 11382 120134
rect 10826 84218 11062 84454
rect 11146 84218 11382 84454
rect 10826 83898 11062 84134
rect 11146 83898 11382 84134
rect 10826 48218 11062 48454
rect 11146 48218 11382 48454
rect 10826 47898 11062 48134
rect 11146 47898 11382 48134
rect 10826 12218 11062 12454
rect 11146 12218 11382 12454
rect 10826 11898 11062 12134
rect 11146 11898 11382 12134
rect 10826 -2502 11062 -2266
rect 11146 -2502 11382 -2266
rect 10826 -2822 11062 -2586
rect 11146 -2822 11382 -2586
rect 15326 707482 15562 707718
rect 15646 707482 15882 707718
rect 15326 707162 15562 707398
rect 15646 707162 15882 707398
rect 15326 700718 15562 700954
rect 15646 700718 15882 700954
rect 15326 700398 15562 700634
rect 15646 700398 15882 700634
rect 15326 664718 15562 664954
rect 15646 664718 15882 664954
rect 15326 664398 15562 664634
rect 15646 664398 15882 664634
rect 15326 628718 15562 628954
rect 15646 628718 15882 628954
rect 15326 628398 15562 628634
rect 15646 628398 15882 628634
rect 15326 592718 15562 592954
rect 15646 592718 15882 592954
rect 15326 592398 15562 592634
rect 15646 592398 15882 592634
rect 15326 556718 15562 556954
rect 15646 556718 15882 556954
rect 15326 556398 15562 556634
rect 15646 556398 15882 556634
rect 15326 520718 15562 520954
rect 15646 520718 15882 520954
rect 15326 520398 15562 520634
rect 15646 520398 15882 520634
rect 15326 484718 15562 484954
rect 15646 484718 15882 484954
rect 15326 484398 15562 484634
rect 15646 484398 15882 484634
rect 15326 448718 15562 448954
rect 15646 448718 15882 448954
rect 15326 448398 15562 448634
rect 15646 448398 15882 448634
rect 15326 412718 15562 412954
rect 15646 412718 15882 412954
rect 15326 412398 15562 412634
rect 15646 412398 15882 412634
rect 15326 376718 15562 376954
rect 15646 376718 15882 376954
rect 15326 376398 15562 376634
rect 15646 376398 15882 376634
rect 15326 340718 15562 340954
rect 15646 340718 15882 340954
rect 15326 340398 15562 340634
rect 15646 340398 15882 340634
rect 15326 304718 15562 304954
rect 15646 304718 15882 304954
rect 15326 304398 15562 304634
rect 15646 304398 15882 304634
rect 15326 268718 15562 268954
rect 15646 268718 15882 268954
rect 15326 268398 15562 268634
rect 15646 268398 15882 268634
rect 15326 232718 15562 232954
rect 15646 232718 15882 232954
rect 15326 232398 15562 232634
rect 15646 232398 15882 232634
rect 15326 196718 15562 196954
rect 15646 196718 15882 196954
rect 15326 196398 15562 196634
rect 15646 196398 15882 196634
rect 15326 160718 15562 160954
rect 15646 160718 15882 160954
rect 15326 160398 15562 160634
rect 15646 160398 15882 160634
rect 15326 124718 15562 124954
rect 15646 124718 15882 124954
rect 15326 124398 15562 124634
rect 15646 124398 15882 124634
rect 15326 88718 15562 88954
rect 15646 88718 15882 88954
rect 15326 88398 15562 88634
rect 15646 88398 15882 88634
rect 15326 52718 15562 52954
rect 15646 52718 15882 52954
rect 15326 52398 15562 52634
rect 15646 52398 15882 52634
rect 15326 16718 15562 16954
rect 15646 16718 15882 16954
rect 15326 16398 15562 16634
rect 15646 16398 15882 16634
rect 15326 -3462 15562 -3226
rect 15646 -3462 15882 -3226
rect 15326 -3782 15562 -3546
rect 15646 -3782 15882 -3546
rect 19826 708442 20062 708678
rect 20146 708442 20382 708678
rect 19826 708122 20062 708358
rect 20146 708122 20382 708358
rect 19826 669218 20062 669454
rect 20146 669218 20382 669454
rect 19826 668898 20062 669134
rect 20146 668898 20382 669134
rect 19826 633218 20062 633454
rect 20146 633218 20382 633454
rect 19826 632898 20062 633134
rect 20146 632898 20382 633134
rect 19826 597218 20062 597454
rect 20146 597218 20382 597454
rect 19826 596898 20062 597134
rect 20146 596898 20382 597134
rect 19826 561218 20062 561454
rect 20146 561218 20382 561454
rect 19826 560898 20062 561134
rect 20146 560898 20382 561134
rect 19826 525218 20062 525454
rect 20146 525218 20382 525454
rect 19826 524898 20062 525134
rect 20146 524898 20382 525134
rect 19826 489218 20062 489454
rect 20146 489218 20382 489454
rect 19826 488898 20062 489134
rect 20146 488898 20382 489134
rect 19826 453218 20062 453454
rect 20146 453218 20382 453454
rect 19826 452898 20062 453134
rect 20146 452898 20382 453134
rect 19826 417218 20062 417454
rect 20146 417218 20382 417454
rect 19826 416898 20062 417134
rect 20146 416898 20382 417134
rect 19826 381218 20062 381454
rect 20146 381218 20382 381454
rect 19826 380898 20062 381134
rect 20146 380898 20382 381134
rect 19826 345218 20062 345454
rect 20146 345218 20382 345454
rect 19826 344898 20062 345134
rect 20146 344898 20382 345134
rect 19826 309218 20062 309454
rect 20146 309218 20382 309454
rect 19826 308898 20062 309134
rect 20146 308898 20382 309134
rect 19826 273218 20062 273454
rect 20146 273218 20382 273454
rect 19826 272898 20062 273134
rect 20146 272898 20382 273134
rect 19826 237218 20062 237454
rect 20146 237218 20382 237454
rect 19826 236898 20062 237134
rect 20146 236898 20382 237134
rect 19826 201218 20062 201454
rect 20146 201218 20382 201454
rect 19826 200898 20062 201134
rect 20146 200898 20382 201134
rect 19826 165218 20062 165454
rect 20146 165218 20382 165454
rect 19826 164898 20062 165134
rect 20146 164898 20382 165134
rect 19826 129218 20062 129454
rect 20146 129218 20382 129454
rect 19826 128898 20062 129134
rect 20146 128898 20382 129134
rect 19826 93218 20062 93454
rect 20146 93218 20382 93454
rect 19826 92898 20062 93134
rect 20146 92898 20382 93134
rect 19826 57218 20062 57454
rect 20146 57218 20382 57454
rect 19826 56898 20062 57134
rect 20146 56898 20382 57134
rect 19826 21218 20062 21454
rect 20146 21218 20382 21454
rect 19826 20898 20062 21134
rect 20146 20898 20382 21134
rect 19826 -4422 20062 -4186
rect 20146 -4422 20382 -4186
rect 19826 -4742 20062 -4506
rect 20146 -4742 20382 -4506
rect 24326 709402 24562 709638
rect 24646 709402 24882 709638
rect 24326 709082 24562 709318
rect 24646 709082 24882 709318
rect 24326 673718 24562 673954
rect 24646 673718 24882 673954
rect 24326 673398 24562 673634
rect 24646 673398 24882 673634
rect 24326 637718 24562 637954
rect 24646 637718 24882 637954
rect 24326 637398 24562 637634
rect 24646 637398 24882 637634
rect 24326 601718 24562 601954
rect 24646 601718 24882 601954
rect 24326 601398 24562 601634
rect 24646 601398 24882 601634
rect 24326 565718 24562 565954
rect 24646 565718 24882 565954
rect 24326 565398 24562 565634
rect 24646 565398 24882 565634
rect 24326 529718 24562 529954
rect 24646 529718 24882 529954
rect 24326 529398 24562 529634
rect 24646 529398 24882 529634
rect 24326 493718 24562 493954
rect 24646 493718 24882 493954
rect 24326 493398 24562 493634
rect 24646 493398 24882 493634
rect 24326 457718 24562 457954
rect 24646 457718 24882 457954
rect 24326 457398 24562 457634
rect 24646 457398 24882 457634
rect 24326 421718 24562 421954
rect 24646 421718 24882 421954
rect 24326 421398 24562 421634
rect 24646 421398 24882 421634
rect 24326 385718 24562 385954
rect 24646 385718 24882 385954
rect 24326 385398 24562 385634
rect 24646 385398 24882 385634
rect 24326 349718 24562 349954
rect 24646 349718 24882 349954
rect 24326 349398 24562 349634
rect 24646 349398 24882 349634
rect 24326 313718 24562 313954
rect 24646 313718 24882 313954
rect 24326 313398 24562 313634
rect 24646 313398 24882 313634
rect 24326 277718 24562 277954
rect 24646 277718 24882 277954
rect 24326 277398 24562 277634
rect 24646 277398 24882 277634
rect 24326 241718 24562 241954
rect 24646 241718 24882 241954
rect 24326 241398 24562 241634
rect 24646 241398 24882 241634
rect 24326 205718 24562 205954
rect 24646 205718 24882 205954
rect 24326 205398 24562 205634
rect 24646 205398 24882 205634
rect 24326 169718 24562 169954
rect 24646 169718 24882 169954
rect 24326 169398 24562 169634
rect 24646 169398 24882 169634
rect 24326 133718 24562 133954
rect 24646 133718 24882 133954
rect 24326 133398 24562 133634
rect 24646 133398 24882 133634
rect 24326 97718 24562 97954
rect 24646 97718 24882 97954
rect 24326 97398 24562 97634
rect 24646 97398 24882 97634
rect 24326 61718 24562 61954
rect 24646 61718 24882 61954
rect 24326 61398 24562 61634
rect 24646 61398 24882 61634
rect 24326 25718 24562 25954
rect 24646 25718 24882 25954
rect 24326 25398 24562 25634
rect 24646 25398 24882 25634
rect 24326 -5382 24562 -5146
rect 24646 -5382 24882 -5146
rect 24326 -5702 24562 -5466
rect 24646 -5702 24882 -5466
rect 28826 710362 29062 710598
rect 29146 710362 29382 710598
rect 28826 710042 29062 710278
rect 29146 710042 29382 710278
rect 28826 678218 29062 678454
rect 29146 678218 29382 678454
rect 28826 677898 29062 678134
rect 29146 677898 29382 678134
rect 28826 642218 29062 642454
rect 29146 642218 29382 642454
rect 28826 641898 29062 642134
rect 29146 641898 29382 642134
rect 28826 606218 29062 606454
rect 29146 606218 29382 606454
rect 28826 605898 29062 606134
rect 29146 605898 29382 606134
rect 28826 570218 29062 570454
rect 29146 570218 29382 570454
rect 28826 569898 29062 570134
rect 29146 569898 29382 570134
rect 28826 534218 29062 534454
rect 29146 534218 29382 534454
rect 28826 533898 29062 534134
rect 29146 533898 29382 534134
rect 28826 498218 29062 498454
rect 29146 498218 29382 498454
rect 28826 497898 29062 498134
rect 29146 497898 29382 498134
rect 28826 462218 29062 462454
rect 29146 462218 29382 462454
rect 28826 461898 29062 462134
rect 29146 461898 29382 462134
rect 28826 426218 29062 426454
rect 29146 426218 29382 426454
rect 28826 425898 29062 426134
rect 29146 425898 29382 426134
rect 28826 390218 29062 390454
rect 29146 390218 29382 390454
rect 28826 389898 29062 390134
rect 29146 389898 29382 390134
rect 28826 354218 29062 354454
rect 29146 354218 29382 354454
rect 28826 353898 29062 354134
rect 29146 353898 29382 354134
rect 28826 318218 29062 318454
rect 29146 318218 29382 318454
rect 28826 317898 29062 318134
rect 29146 317898 29382 318134
rect 28826 282218 29062 282454
rect 29146 282218 29382 282454
rect 28826 281898 29062 282134
rect 29146 281898 29382 282134
rect 28826 246218 29062 246454
rect 29146 246218 29382 246454
rect 28826 245898 29062 246134
rect 29146 245898 29382 246134
rect 28826 210218 29062 210454
rect 29146 210218 29382 210454
rect 28826 209898 29062 210134
rect 29146 209898 29382 210134
rect 28826 174218 29062 174454
rect 29146 174218 29382 174454
rect 28826 173898 29062 174134
rect 29146 173898 29382 174134
rect 28826 138218 29062 138454
rect 29146 138218 29382 138454
rect 28826 137898 29062 138134
rect 29146 137898 29382 138134
rect 28826 102218 29062 102454
rect 29146 102218 29382 102454
rect 28826 101898 29062 102134
rect 29146 101898 29382 102134
rect 28826 66218 29062 66454
rect 29146 66218 29382 66454
rect 28826 65898 29062 66134
rect 29146 65898 29382 66134
rect 28826 30218 29062 30454
rect 29146 30218 29382 30454
rect 28826 29898 29062 30134
rect 29146 29898 29382 30134
rect 28826 -6342 29062 -6106
rect 29146 -6342 29382 -6106
rect 28826 -6662 29062 -6426
rect 29146 -6662 29382 -6426
rect 33326 711322 33562 711558
rect 33646 711322 33882 711558
rect 33326 711002 33562 711238
rect 33646 711002 33882 711238
rect 33326 682718 33562 682954
rect 33646 682718 33882 682954
rect 33326 682398 33562 682634
rect 33646 682398 33882 682634
rect 33326 646718 33562 646954
rect 33646 646718 33882 646954
rect 33326 646398 33562 646634
rect 33646 646398 33882 646634
rect 33326 610718 33562 610954
rect 33646 610718 33882 610954
rect 33326 610398 33562 610634
rect 33646 610398 33882 610634
rect 33326 574718 33562 574954
rect 33646 574718 33882 574954
rect 33326 574398 33562 574634
rect 33646 574398 33882 574634
rect 33326 538718 33562 538954
rect 33646 538718 33882 538954
rect 33326 538398 33562 538634
rect 33646 538398 33882 538634
rect 33326 502718 33562 502954
rect 33646 502718 33882 502954
rect 33326 502398 33562 502634
rect 33646 502398 33882 502634
rect 33326 466718 33562 466954
rect 33646 466718 33882 466954
rect 33326 466398 33562 466634
rect 33646 466398 33882 466634
rect 33326 430718 33562 430954
rect 33646 430718 33882 430954
rect 33326 430398 33562 430634
rect 33646 430398 33882 430634
rect 33326 394718 33562 394954
rect 33646 394718 33882 394954
rect 33326 394398 33562 394634
rect 33646 394398 33882 394634
rect 33326 358718 33562 358954
rect 33646 358718 33882 358954
rect 33326 358398 33562 358634
rect 33646 358398 33882 358634
rect 33326 322718 33562 322954
rect 33646 322718 33882 322954
rect 33326 322398 33562 322634
rect 33646 322398 33882 322634
rect 33326 286718 33562 286954
rect 33646 286718 33882 286954
rect 33326 286398 33562 286634
rect 33646 286398 33882 286634
rect 33326 250718 33562 250954
rect 33646 250718 33882 250954
rect 33326 250398 33562 250634
rect 33646 250398 33882 250634
rect 33326 214718 33562 214954
rect 33646 214718 33882 214954
rect 33326 214398 33562 214634
rect 33646 214398 33882 214634
rect 33326 178718 33562 178954
rect 33646 178718 33882 178954
rect 33326 178398 33562 178634
rect 33646 178398 33882 178634
rect 33326 142718 33562 142954
rect 33646 142718 33882 142954
rect 33326 142398 33562 142634
rect 33646 142398 33882 142634
rect 33326 106718 33562 106954
rect 33646 106718 33882 106954
rect 33326 106398 33562 106634
rect 33646 106398 33882 106634
rect 33326 70718 33562 70954
rect 33646 70718 33882 70954
rect 33326 70398 33562 70634
rect 33646 70398 33882 70634
rect 33326 34718 33562 34954
rect 33646 34718 33882 34954
rect 33326 34398 33562 34634
rect 33646 34398 33882 34634
rect 33326 -7302 33562 -7066
rect 33646 -7302 33882 -7066
rect 33326 -7622 33562 -7386
rect 33646 -7622 33882 -7386
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 37826 651218 38062 651454
rect 38146 651218 38382 651454
rect 37826 650898 38062 651134
rect 38146 650898 38382 651134
rect 37826 615218 38062 615454
rect 38146 615218 38382 615454
rect 37826 614898 38062 615134
rect 38146 614898 38382 615134
rect 37826 579218 38062 579454
rect 38146 579218 38382 579454
rect 37826 578898 38062 579134
rect 38146 578898 38382 579134
rect 37826 543218 38062 543454
rect 38146 543218 38382 543454
rect 37826 542898 38062 543134
rect 38146 542898 38382 543134
rect 37826 507218 38062 507454
rect 38146 507218 38382 507454
rect 37826 506898 38062 507134
rect 38146 506898 38382 507134
rect 37826 471218 38062 471454
rect 38146 471218 38382 471454
rect 37826 470898 38062 471134
rect 38146 470898 38382 471134
rect 37826 435218 38062 435454
rect 38146 435218 38382 435454
rect 37826 434898 38062 435134
rect 38146 434898 38382 435134
rect 37826 399218 38062 399454
rect 38146 399218 38382 399454
rect 37826 398898 38062 399134
rect 38146 398898 38382 399134
rect 37826 363218 38062 363454
rect 38146 363218 38382 363454
rect 37826 362898 38062 363134
rect 38146 362898 38382 363134
rect 37826 327218 38062 327454
rect 38146 327218 38382 327454
rect 37826 326898 38062 327134
rect 38146 326898 38382 327134
rect 37826 291218 38062 291454
rect 38146 291218 38382 291454
rect 37826 290898 38062 291134
rect 38146 290898 38382 291134
rect 37826 255218 38062 255454
rect 38146 255218 38382 255454
rect 37826 254898 38062 255134
rect 38146 254898 38382 255134
rect 37826 219218 38062 219454
rect 38146 219218 38382 219454
rect 37826 218898 38062 219134
rect 38146 218898 38382 219134
rect 37826 183218 38062 183454
rect 38146 183218 38382 183454
rect 37826 182898 38062 183134
rect 38146 182898 38382 183134
rect 37826 147218 38062 147454
rect 38146 147218 38382 147454
rect 37826 146898 38062 147134
rect 38146 146898 38382 147134
rect 37826 111218 38062 111454
rect 38146 111218 38382 111454
rect 37826 110898 38062 111134
rect 38146 110898 38382 111134
rect 37826 75218 38062 75454
rect 38146 75218 38382 75454
rect 37826 74898 38062 75134
rect 38146 74898 38382 75134
rect 37826 39218 38062 39454
rect 38146 39218 38382 39454
rect 37826 38898 38062 39134
rect 38146 38898 38382 39134
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 42326 705562 42562 705798
rect 42646 705562 42882 705798
rect 42326 705242 42562 705478
rect 42646 705242 42882 705478
rect 42326 691718 42562 691954
rect 42646 691718 42882 691954
rect 42326 691398 42562 691634
rect 42646 691398 42882 691634
rect 42326 655718 42562 655954
rect 42646 655718 42882 655954
rect 42326 655398 42562 655634
rect 42646 655398 42882 655634
rect 42326 619718 42562 619954
rect 42646 619718 42882 619954
rect 42326 619398 42562 619634
rect 42646 619398 42882 619634
rect 42326 583718 42562 583954
rect 42646 583718 42882 583954
rect 42326 583398 42562 583634
rect 42646 583398 42882 583634
rect 42326 547718 42562 547954
rect 42646 547718 42882 547954
rect 42326 547398 42562 547634
rect 42646 547398 42882 547634
rect 42326 511718 42562 511954
rect 42646 511718 42882 511954
rect 42326 511398 42562 511634
rect 42646 511398 42882 511634
rect 42326 475718 42562 475954
rect 42646 475718 42882 475954
rect 42326 475398 42562 475634
rect 42646 475398 42882 475634
rect 42326 439718 42562 439954
rect 42646 439718 42882 439954
rect 42326 439398 42562 439634
rect 42646 439398 42882 439634
rect 42326 403718 42562 403954
rect 42646 403718 42882 403954
rect 42326 403398 42562 403634
rect 42646 403398 42882 403634
rect 42326 367718 42562 367954
rect 42646 367718 42882 367954
rect 42326 367398 42562 367634
rect 42646 367398 42882 367634
rect 42326 331718 42562 331954
rect 42646 331718 42882 331954
rect 42326 331398 42562 331634
rect 42646 331398 42882 331634
rect 42326 295718 42562 295954
rect 42646 295718 42882 295954
rect 42326 295398 42562 295634
rect 42646 295398 42882 295634
rect 42326 259718 42562 259954
rect 42646 259718 42882 259954
rect 42326 259398 42562 259634
rect 42646 259398 42882 259634
rect 42326 223718 42562 223954
rect 42646 223718 42882 223954
rect 42326 223398 42562 223634
rect 42646 223398 42882 223634
rect 42326 187718 42562 187954
rect 42646 187718 42882 187954
rect 42326 187398 42562 187634
rect 42646 187398 42882 187634
rect 42326 151718 42562 151954
rect 42646 151718 42882 151954
rect 42326 151398 42562 151634
rect 42646 151398 42882 151634
rect 42326 115718 42562 115954
rect 42646 115718 42882 115954
rect 42326 115398 42562 115634
rect 42646 115398 42882 115634
rect 42326 79718 42562 79954
rect 42646 79718 42882 79954
rect 42326 79398 42562 79634
rect 42646 79398 42882 79634
rect 42326 43718 42562 43954
rect 42646 43718 42882 43954
rect 42326 43398 42562 43634
rect 42646 43398 42882 43634
rect 42326 7718 42562 7954
rect 42646 7718 42882 7954
rect 42326 7398 42562 7634
rect 42646 7398 42882 7634
rect 42326 -1542 42562 -1306
rect 42646 -1542 42882 -1306
rect 42326 -1862 42562 -1626
rect 42646 -1862 42882 -1626
rect 46826 706522 47062 706758
rect 47146 706522 47382 706758
rect 46826 706202 47062 706438
rect 47146 706202 47382 706438
rect 46826 696218 47062 696454
rect 47146 696218 47382 696454
rect 46826 695898 47062 696134
rect 47146 695898 47382 696134
rect 46826 660218 47062 660454
rect 47146 660218 47382 660454
rect 46826 659898 47062 660134
rect 47146 659898 47382 660134
rect 46826 624218 47062 624454
rect 47146 624218 47382 624454
rect 46826 623898 47062 624134
rect 47146 623898 47382 624134
rect 46826 588218 47062 588454
rect 47146 588218 47382 588454
rect 46826 587898 47062 588134
rect 47146 587898 47382 588134
rect 46826 552218 47062 552454
rect 47146 552218 47382 552454
rect 46826 551898 47062 552134
rect 47146 551898 47382 552134
rect 46826 516218 47062 516454
rect 47146 516218 47382 516454
rect 46826 515898 47062 516134
rect 47146 515898 47382 516134
rect 46826 480218 47062 480454
rect 47146 480218 47382 480454
rect 46826 479898 47062 480134
rect 47146 479898 47382 480134
rect 46826 444218 47062 444454
rect 47146 444218 47382 444454
rect 46826 443898 47062 444134
rect 47146 443898 47382 444134
rect 46826 408218 47062 408454
rect 47146 408218 47382 408454
rect 46826 407898 47062 408134
rect 47146 407898 47382 408134
rect 46826 372218 47062 372454
rect 47146 372218 47382 372454
rect 46826 371898 47062 372134
rect 47146 371898 47382 372134
rect 46826 336218 47062 336454
rect 47146 336218 47382 336454
rect 46826 335898 47062 336134
rect 47146 335898 47382 336134
rect 46826 300218 47062 300454
rect 47146 300218 47382 300454
rect 46826 299898 47062 300134
rect 47146 299898 47382 300134
rect 46826 264218 47062 264454
rect 47146 264218 47382 264454
rect 46826 263898 47062 264134
rect 47146 263898 47382 264134
rect 46826 228218 47062 228454
rect 47146 228218 47382 228454
rect 46826 227898 47062 228134
rect 47146 227898 47382 228134
rect 46826 192218 47062 192454
rect 47146 192218 47382 192454
rect 46826 191898 47062 192134
rect 47146 191898 47382 192134
rect 46826 156218 47062 156454
rect 47146 156218 47382 156454
rect 46826 155898 47062 156134
rect 47146 155898 47382 156134
rect 46826 120218 47062 120454
rect 47146 120218 47382 120454
rect 46826 119898 47062 120134
rect 47146 119898 47382 120134
rect 46826 84218 47062 84454
rect 47146 84218 47382 84454
rect 46826 83898 47062 84134
rect 47146 83898 47382 84134
rect 46826 48218 47062 48454
rect 47146 48218 47382 48454
rect 46826 47898 47062 48134
rect 47146 47898 47382 48134
rect 46826 12218 47062 12454
rect 47146 12218 47382 12454
rect 46826 11898 47062 12134
rect 47146 11898 47382 12134
rect 46826 -2502 47062 -2266
rect 47146 -2502 47382 -2266
rect 46826 -2822 47062 -2586
rect 47146 -2822 47382 -2586
rect 51326 707482 51562 707718
rect 51646 707482 51882 707718
rect 51326 707162 51562 707398
rect 51646 707162 51882 707398
rect 51326 700718 51562 700954
rect 51646 700718 51882 700954
rect 51326 700398 51562 700634
rect 51646 700398 51882 700634
rect 51326 664718 51562 664954
rect 51646 664718 51882 664954
rect 51326 664398 51562 664634
rect 51646 664398 51882 664634
rect 51326 628718 51562 628954
rect 51646 628718 51882 628954
rect 51326 628398 51562 628634
rect 51646 628398 51882 628634
rect 51326 592718 51562 592954
rect 51646 592718 51882 592954
rect 51326 592398 51562 592634
rect 51646 592398 51882 592634
rect 51326 556718 51562 556954
rect 51646 556718 51882 556954
rect 51326 556398 51562 556634
rect 51646 556398 51882 556634
rect 51326 520718 51562 520954
rect 51646 520718 51882 520954
rect 51326 520398 51562 520634
rect 51646 520398 51882 520634
rect 51326 484718 51562 484954
rect 51646 484718 51882 484954
rect 51326 484398 51562 484634
rect 51646 484398 51882 484634
rect 51326 448718 51562 448954
rect 51646 448718 51882 448954
rect 51326 448398 51562 448634
rect 51646 448398 51882 448634
rect 51326 412718 51562 412954
rect 51646 412718 51882 412954
rect 51326 412398 51562 412634
rect 51646 412398 51882 412634
rect 51326 376718 51562 376954
rect 51646 376718 51882 376954
rect 51326 376398 51562 376634
rect 51646 376398 51882 376634
rect 51326 340718 51562 340954
rect 51646 340718 51882 340954
rect 51326 340398 51562 340634
rect 51646 340398 51882 340634
rect 51326 304718 51562 304954
rect 51646 304718 51882 304954
rect 51326 304398 51562 304634
rect 51646 304398 51882 304634
rect 51326 268718 51562 268954
rect 51646 268718 51882 268954
rect 51326 268398 51562 268634
rect 51646 268398 51882 268634
rect 51326 232718 51562 232954
rect 51646 232718 51882 232954
rect 51326 232398 51562 232634
rect 51646 232398 51882 232634
rect 51326 196718 51562 196954
rect 51646 196718 51882 196954
rect 51326 196398 51562 196634
rect 51646 196398 51882 196634
rect 51326 160718 51562 160954
rect 51646 160718 51882 160954
rect 51326 160398 51562 160634
rect 51646 160398 51882 160634
rect 51326 124718 51562 124954
rect 51646 124718 51882 124954
rect 51326 124398 51562 124634
rect 51646 124398 51882 124634
rect 51326 88718 51562 88954
rect 51646 88718 51882 88954
rect 51326 88398 51562 88634
rect 51646 88398 51882 88634
rect 51326 52718 51562 52954
rect 51646 52718 51882 52954
rect 51326 52398 51562 52634
rect 51646 52398 51882 52634
rect 51326 16718 51562 16954
rect 51646 16718 51882 16954
rect 51326 16398 51562 16634
rect 51646 16398 51882 16634
rect 51326 -3462 51562 -3226
rect 51646 -3462 51882 -3226
rect 51326 -3782 51562 -3546
rect 51646 -3782 51882 -3546
rect 55826 708442 56062 708678
rect 56146 708442 56382 708678
rect 55826 708122 56062 708358
rect 56146 708122 56382 708358
rect 55826 669218 56062 669454
rect 56146 669218 56382 669454
rect 55826 668898 56062 669134
rect 56146 668898 56382 669134
rect 55826 633218 56062 633454
rect 56146 633218 56382 633454
rect 55826 632898 56062 633134
rect 56146 632898 56382 633134
rect 55826 597218 56062 597454
rect 56146 597218 56382 597454
rect 55826 596898 56062 597134
rect 56146 596898 56382 597134
rect 55826 561218 56062 561454
rect 56146 561218 56382 561454
rect 55826 560898 56062 561134
rect 56146 560898 56382 561134
rect 55826 525218 56062 525454
rect 56146 525218 56382 525454
rect 55826 524898 56062 525134
rect 56146 524898 56382 525134
rect 55826 489218 56062 489454
rect 56146 489218 56382 489454
rect 55826 488898 56062 489134
rect 56146 488898 56382 489134
rect 55826 453218 56062 453454
rect 56146 453218 56382 453454
rect 55826 452898 56062 453134
rect 56146 452898 56382 453134
rect 55826 417218 56062 417454
rect 56146 417218 56382 417454
rect 55826 416898 56062 417134
rect 56146 416898 56382 417134
rect 55826 381218 56062 381454
rect 56146 381218 56382 381454
rect 55826 380898 56062 381134
rect 56146 380898 56382 381134
rect 55826 345218 56062 345454
rect 56146 345218 56382 345454
rect 55826 344898 56062 345134
rect 56146 344898 56382 345134
rect 55826 309218 56062 309454
rect 56146 309218 56382 309454
rect 55826 308898 56062 309134
rect 56146 308898 56382 309134
rect 55826 273218 56062 273454
rect 56146 273218 56382 273454
rect 55826 272898 56062 273134
rect 56146 272898 56382 273134
rect 55826 237218 56062 237454
rect 56146 237218 56382 237454
rect 55826 236898 56062 237134
rect 56146 236898 56382 237134
rect 55826 201218 56062 201454
rect 56146 201218 56382 201454
rect 55826 200898 56062 201134
rect 56146 200898 56382 201134
rect 55826 165218 56062 165454
rect 56146 165218 56382 165454
rect 55826 164898 56062 165134
rect 56146 164898 56382 165134
rect 55826 129218 56062 129454
rect 56146 129218 56382 129454
rect 55826 128898 56062 129134
rect 56146 128898 56382 129134
rect 55826 93218 56062 93454
rect 56146 93218 56382 93454
rect 55826 92898 56062 93134
rect 56146 92898 56382 93134
rect 55826 57218 56062 57454
rect 56146 57218 56382 57454
rect 55826 56898 56062 57134
rect 56146 56898 56382 57134
rect 55826 21218 56062 21454
rect 56146 21218 56382 21454
rect 55826 20898 56062 21134
rect 56146 20898 56382 21134
rect 55826 -4422 56062 -4186
rect 56146 -4422 56382 -4186
rect 55826 -4742 56062 -4506
rect 56146 -4742 56382 -4506
rect 60326 709402 60562 709638
rect 60646 709402 60882 709638
rect 60326 709082 60562 709318
rect 60646 709082 60882 709318
rect 60326 673718 60562 673954
rect 60646 673718 60882 673954
rect 60326 673398 60562 673634
rect 60646 673398 60882 673634
rect 60326 637718 60562 637954
rect 60646 637718 60882 637954
rect 60326 637398 60562 637634
rect 60646 637398 60882 637634
rect 60326 601718 60562 601954
rect 60646 601718 60882 601954
rect 60326 601398 60562 601634
rect 60646 601398 60882 601634
rect 60326 565718 60562 565954
rect 60646 565718 60882 565954
rect 60326 565398 60562 565634
rect 60646 565398 60882 565634
rect 60326 529718 60562 529954
rect 60646 529718 60882 529954
rect 60326 529398 60562 529634
rect 60646 529398 60882 529634
rect 60326 493718 60562 493954
rect 60646 493718 60882 493954
rect 60326 493398 60562 493634
rect 60646 493398 60882 493634
rect 60326 457718 60562 457954
rect 60646 457718 60882 457954
rect 60326 457398 60562 457634
rect 60646 457398 60882 457634
rect 60326 421718 60562 421954
rect 60646 421718 60882 421954
rect 60326 421398 60562 421634
rect 60646 421398 60882 421634
rect 60326 385718 60562 385954
rect 60646 385718 60882 385954
rect 60326 385398 60562 385634
rect 60646 385398 60882 385634
rect 60326 349718 60562 349954
rect 60646 349718 60882 349954
rect 60326 349398 60562 349634
rect 60646 349398 60882 349634
rect 60326 313718 60562 313954
rect 60646 313718 60882 313954
rect 60326 313398 60562 313634
rect 60646 313398 60882 313634
rect 60326 277718 60562 277954
rect 60646 277718 60882 277954
rect 60326 277398 60562 277634
rect 60646 277398 60882 277634
rect 60326 241718 60562 241954
rect 60646 241718 60882 241954
rect 60326 241398 60562 241634
rect 60646 241398 60882 241634
rect 60326 205718 60562 205954
rect 60646 205718 60882 205954
rect 60326 205398 60562 205634
rect 60646 205398 60882 205634
rect 60326 169718 60562 169954
rect 60646 169718 60882 169954
rect 60326 169398 60562 169634
rect 60646 169398 60882 169634
rect 60326 133718 60562 133954
rect 60646 133718 60882 133954
rect 60326 133398 60562 133634
rect 60646 133398 60882 133634
rect 60326 97718 60562 97954
rect 60646 97718 60882 97954
rect 60326 97398 60562 97634
rect 60646 97398 60882 97634
rect 60326 61718 60562 61954
rect 60646 61718 60882 61954
rect 60326 61398 60562 61634
rect 60646 61398 60882 61634
rect 60326 25718 60562 25954
rect 60646 25718 60882 25954
rect 60326 25398 60562 25634
rect 60646 25398 60882 25634
rect 60326 -5382 60562 -5146
rect 60646 -5382 60882 -5146
rect 60326 -5702 60562 -5466
rect 60646 -5702 60882 -5466
rect 64826 710362 65062 710598
rect 65146 710362 65382 710598
rect 64826 710042 65062 710278
rect 65146 710042 65382 710278
rect 64826 678218 65062 678454
rect 65146 678218 65382 678454
rect 64826 677898 65062 678134
rect 65146 677898 65382 678134
rect 64826 642218 65062 642454
rect 65146 642218 65382 642454
rect 64826 641898 65062 642134
rect 65146 641898 65382 642134
rect 64826 606218 65062 606454
rect 65146 606218 65382 606454
rect 64826 605898 65062 606134
rect 65146 605898 65382 606134
rect 64826 570218 65062 570454
rect 65146 570218 65382 570454
rect 64826 569898 65062 570134
rect 65146 569898 65382 570134
rect 64826 534218 65062 534454
rect 65146 534218 65382 534454
rect 64826 533898 65062 534134
rect 65146 533898 65382 534134
rect 64826 498218 65062 498454
rect 65146 498218 65382 498454
rect 64826 497898 65062 498134
rect 65146 497898 65382 498134
rect 64826 462218 65062 462454
rect 65146 462218 65382 462454
rect 64826 461898 65062 462134
rect 65146 461898 65382 462134
rect 64826 426218 65062 426454
rect 65146 426218 65382 426454
rect 64826 425898 65062 426134
rect 65146 425898 65382 426134
rect 64826 390218 65062 390454
rect 65146 390218 65382 390454
rect 64826 389898 65062 390134
rect 65146 389898 65382 390134
rect 64826 354218 65062 354454
rect 65146 354218 65382 354454
rect 64826 353898 65062 354134
rect 65146 353898 65382 354134
rect 64826 318218 65062 318454
rect 65146 318218 65382 318454
rect 64826 317898 65062 318134
rect 65146 317898 65382 318134
rect 64826 282218 65062 282454
rect 65146 282218 65382 282454
rect 64826 281898 65062 282134
rect 65146 281898 65382 282134
rect 64826 246218 65062 246454
rect 65146 246218 65382 246454
rect 64826 245898 65062 246134
rect 65146 245898 65382 246134
rect 64826 210218 65062 210454
rect 65146 210218 65382 210454
rect 64826 209898 65062 210134
rect 65146 209898 65382 210134
rect 64826 174218 65062 174454
rect 65146 174218 65382 174454
rect 64826 173898 65062 174134
rect 65146 173898 65382 174134
rect 64826 138218 65062 138454
rect 65146 138218 65382 138454
rect 64826 137898 65062 138134
rect 65146 137898 65382 138134
rect 64826 102218 65062 102454
rect 65146 102218 65382 102454
rect 64826 101898 65062 102134
rect 65146 101898 65382 102134
rect 64826 66218 65062 66454
rect 65146 66218 65382 66454
rect 64826 65898 65062 66134
rect 65146 65898 65382 66134
rect 64826 30218 65062 30454
rect 65146 30218 65382 30454
rect 64826 29898 65062 30134
rect 65146 29898 65382 30134
rect 64826 -6342 65062 -6106
rect 65146 -6342 65382 -6106
rect 64826 -6662 65062 -6426
rect 65146 -6662 65382 -6426
rect 69326 711322 69562 711558
rect 69646 711322 69882 711558
rect 69326 711002 69562 711238
rect 69646 711002 69882 711238
rect 69326 682718 69562 682954
rect 69646 682718 69882 682954
rect 69326 682398 69562 682634
rect 69646 682398 69882 682634
rect 69326 646718 69562 646954
rect 69646 646718 69882 646954
rect 69326 646398 69562 646634
rect 69646 646398 69882 646634
rect 69326 610718 69562 610954
rect 69646 610718 69882 610954
rect 69326 610398 69562 610634
rect 69646 610398 69882 610634
rect 69326 574718 69562 574954
rect 69646 574718 69882 574954
rect 69326 574398 69562 574634
rect 69646 574398 69882 574634
rect 69326 538718 69562 538954
rect 69646 538718 69882 538954
rect 69326 538398 69562 538634
rect 69646 538398 69882 538634
rect 69326 502718 69562 502954
rect 69646 502718 69882 502954
rect 69326 502398 69562 502634
rect 69646 502398 69882 502634
rect 69326 466718 69562 466954
rect 69646 466718 69882 466954
rect 69326 466398 69562 466634
rect 69646 466398 69882 466634
rect 69326 430718 69562 430954
rect 69646 430718 69882 430954
rect 69326 430398 69562 430634
rect 69646 430398 69882 430634
rect 69326 394718 69562 394954
rect 69646 394718 69882 394954
rect 69326 394398 69562 394634
rect 69646 394398 69882 394634
rect 69326 358718 69562 358954
rect 69646 358718 69882 358954
rect 69326 358398 69562 358634
rect 69646 358398 69882 358634
rect 69326 322718 69562 322954
rect 69646 322718 69882 322954
rect 69326 322398 69562 322634
rect 69646 322398 69882 322634
rect 69326 286718 69562 286954
rect 69646 286718 69882 286954
rect 69326 286398 69562 286634
rect 69646 286398 69882 286634
rect 69326 250718 69562 250954
rect 69646 250718 69882 250954
rect 69326 250398 69562 250634
rect 69646 250398 69882 250634
rect 69326 214718 69562 214954
rect 69646 214718 69882 214954
rect 69326 214398 69562 214634
rect 69646 214398 69882 214634
rect 69326 178718 69562 178954
rect 69646 178718 69882 178954
rect 69326 178398 69562 178634
rect 69646 178398 69882 178634
rect 69326 142718 69562 142954
rect 69646 142718 69882 142954
rect 69326 142398 69562 142634
rect 69646 142398 69882 142634
rect 69326 106718 69562 106954
rect 69646 106718 69882 106954
rect 69326 106398 69562 106634
rect 69646 106398 69882 106634
rect 69326 70718 69562 70954
rect 69646 70718 69882 70954
rect 69326 70398 69562 70634
rect 69646 70398 69882 70634
rect 69326 34718 69562 34954
rect 69646 34718 69882 34954
rect 69326 34398 69562 34634
rect 69646 34398 69882 34634
rect 69326 -7302 69562 -7066
rect 69646 -7302 69882 -7066
rect 69326 -7622 69562 -7386
rect 69646 -7622 69882 -7386
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 73826 651218 74062 651454
rect 74146 651218 74382 651454
rect 73826 650898 74062 651134
rect 74146 650898 74382 651134
rect 73826 615218 74062 615454
rect 74146 615218 74382 615454
rect 73826 614898 74062 615134
rect 74146 614898 74382 615134
rect 73826 579218 74062 579454
rect 74146 579218 74382 579454
rect 73826 578898 74062 579134
rect 74146 578898 74382 579134
rect 73826 543218 74062 543454
rect 74146 543218 74382 543454
rect 73826 542898 74062 543134
rect 74146 542898 74382 543134
rect 73826 507218 74062 507454
rect 74146 507218 74382 507454
rect 73826 506898 74062 507134
rect 74146 506898 74382 507134
rect 73826 471218 74062 471454
rect 74146 471218 74382 471454
rect 73826 470898 74062 471134
rect 74146 470898 74382 471134
rect 73826 435218 74062 435454
rect 74146 435218 74382 435454
rect 73826 434898 74062 435134
rect 74146 434898 74382 435134
rect 73826 399218 74062 399454
rect 74146 399218 74382 399454
rect 73826 398898 74062 399134
rect 74146 398898 74382 399134
rect 73826 363218 74062 363454
rect 74146 363218 74382 363454
rect 73826 362898 74062 363134
rect 74146 362898 74382 363134
rect 73826 327218 74062 327454
rect 74146 327218 74382 327454
rect 73826 326898 74062 327134
rect 74146 326898 74382 327134
rect 73826 291218 74062 291454
rect 74146 291218 74382 291454
rect 73826 290898 74062 291134
rect 74146 290898 74382 291134
rect 73826 255218 74062 255454
rect 74146 255218 74382 255454
rect 73826 254898 74062 255134
rect 74146 254898 74382 255134
rect 73826 219218 74062 219454
rect 74146 219218 74382 219454
rect 73826 218898 74062 219134
rect 74146 218898 74382 219134
rect 73826 183218 74062 183454
rect 74146 183218 74382 183454
rect 73826 182898 74062 183134
rect 74146 182898 74382 183134
rect 73826 147218 74062 147454
rect 74146 147218 74382 147454
rect 73826 146898 74062 147134
rect 74146 146898 74382 147134
rect 73826 111218 74062 111454
rect 74146 111218 74382 111454
rect 73826 110898 74062 111134
rect 74146 110898 74382 111134
rect 73826 75218 74062 75454
rect 74146 75218 74382 75454
rect 73826 74898 74062 75134
rect 74146 74898 74382 75134
rect 73826 39218 74062 39454
rect 74146 39218 74382 39454
rect 73826 38898 74062 39134
rect 74146 38898 74382 39134
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 78326 705562 78562 705798
rect 78646 705562 78882 705798
rect 78326 705242 78562 705478
rect 78646 705242 78882 705478
rect 78326 691718 78562 691954
rect 78646 691718 78882 691954
rect 78326 691398 78562 691634
rect 78646 691398 78882 691634
rect 78326 655718 78562 655954
rect 78646 655718 78882 655954
rect 78326 655398 78562 655634
rect 78646 655398 78882 655634
rect 78326 619718 78562 619954
rect 78646 619718 78882 619954
rect 78326 619398 78562 619634
rect 78646 619398 78882 619634
rect 78326 583718 78562 583954
rect 78646 583718 78882 583954
rect 78326 583398 78562 583634
rect 78646 583398 78882 583634
rect 78326 547718 78562 547954
rect 78646 547718 78882 547954
rect 78326 547398 78562 547634
rect 78646 547398 78882 547634
rect 78326 511718 78562 511954
rect 78646 511718 78882 511954
rect 78326 511398 78562 511634
rect 78646 511398 78882 511634
rect 78326 475718 78562 475954
rect 78646 475718 78882 475954
rect 78326 475398 78562 475634
rect 78646 475398 78882 475634
rect 78326 439718 78562 439954
rect 78646 439718 78882 439954
rect 78326 439398 78562 439634
rect 78646 439398 78882 439634
rect 78326 403718 78562 403954
rect 78646 403718 78882 403954
rect 78326 403398 78562 403634
rect 78646 403398 78882 403634
rect 78326 367718 78562 367954
rect 78646 367718 78882 367954
rect 78326 367398 78562 367634
rect 78646 367398 78882 367634
rect 78326 331718 78562 331954
rect 78646 331718 78882 331954
rect 78326 331398 78562 331634
rect 78646 331398 78882 331634
rect 78326 295718 78562 295954
rect 78646 295718 78882 295954
rect 78326 295398 78562 295634
rect 78646 295398 78882 295634
rect 78326 259718 78562 259954
rect 78646 259718 78882 259954
rect 78326 259398 78562 259634
rect 78646 259398 78882 259634
rect 78326 223718 78562 223954
rect 78646 223718 78882 223954
rect 78326 223398 78562 223634
rect 78646 223398 78882 223634
rect 78326 187718 78562 187954
rect 78646 187718 78882 187954
rect 78326 187398 78562 187634
rect 78646 187398 78882 187634
rect 78326 151718 78562 151954
rect 78646 151718 78882 151954
rect 78326 151398 78562 151634
rect 78646 151398 78882 151634
rect 78326 115718 78562 115954
rect 78646 115718 78882 115954
rect 78326 115398 78562 115634
rect 78646 115398 78882 115634
rect 78326 79718 78562 79954
rect 78646 79718 78882 79954
rect 78326 79398 78562 79634
rect 78646 79398 78882 79634
rect 78326 43718 78562 43954
rect 78646 43718 78882 43954
rect 78326 43398 78562 43634
rect 78646 43398 78882 43634
rect 78326 7718 78562 7954
rect 78646 7718 78882 7954
rect 78326 7398 78562 7634
rect 78646 7398 78882 7634
rect 78326 -1542 78562 -1306
rect 78646 -1542 78882 -1306
rect 78326 -1862 78562 -1626
rect 78646 -1862 78882 -1626
rect 82826 706522 83062 706758
rect 83146 706522 83382 706758
rect 82826 706202 83062 706438
rect 83146 706202 83382 706438
rect 82826 696218 83062 696454
rect 83146 696218 83382 696454
rect 82826 695898 83062 696134
rect 83146 695898 83382 696134
rect 82826 660218 83062 660454
rect 83146 660218 83382 660454
rect 82826 659898 83062 660134
rect 83146 659898 83382 660134
rect 82826 624218 83062 624454
rect 83146 624218 83382 624454
rect 82826 623898 83062 624134
rect 83146 623898 83382 624134
rect 82826 588218 83062 588454
rect 83146 588218 83382 588454
rect 82826 587898 83062 588134
rect 83146 587898 83382 588134
rect 82826 552218 83062 552454
rect 83146 552218 83382 552454
rect 82826 551898 83062 552134
rect 83146 551898 83382 552134
rect 82826 516218 83062 516454
rect 83146 516218 83382 516454
rect 82826 515898 83062 516134
rect 83146 515898 83382 516134
rect 82826 480218 83062 480454
rect 83146 480218 83382 480454
rect 82826 479898 83062 480134
rect 83146 479898 83382 480134
rect 82826 444218 83062 444454
rect 83146 444218 83382 444454
rect 82826 443898 83062 444134
rect 83146 443898 83382 444134
rect 82826 408218 83062 408454
rect 83146 408218 83382 408454
rect 82826 407898 83062 408134
rect 83146 407898 83382 408134
rect 82826 372218 83062 372454
rect 83146 372218 83382 372454
rect 82826 371898 83062 372134
rect 83146 371898 83382 372134
rect 82826 336218 83062 336454
rect 83146 336218 83382 336454
rect 82826 335898 83062 336134
rect 83146 335898 83382 336134
rect 82826 300218 83062 300454
rect 83146 300218 83382 300454
rect 82826 299898 83062 300134
rect 83146 299898 83382 300134
rect 82826 264218 83062 264454
rect 83146 264218 83382 264454
rect 82826 263898 83062 264134
rect 83146 263898 83382 264134
rect 82826 228218 83062 228454
rect 83146 228218 83382 228454
rect 82826 227898 83062 228134
rect 83146 227898 83382 228134
rect 82826 192218 83062 192454
rect 83146 192218 83382 192454
rect 82826 191898 83062 192134
rect 83146 191898 83382 192134
rect 82826 156218 83062 156454
rect 83146 156218 83382 156454
rect 82826 155898 83062 156134
rect 83146 155898 83382 156134
rect 82826 120218 83062 120454
rect 83146 120218 83382 120454
rect 82826 119898 83062 120134
rect 83146 119898 83382 120134
rect 82826 84218 83062 84454
rect 83146 84218 83382 84454
rect 82826 83898 83062 84134
rect 83146 83898 83382 84134
rect 82826 48218 83062 48454
rect 83146 48218 83382 48454
rect 82826 47898 83062 48134
rect 83146 47898 83382 48134
rect 82826 12218 83062 12454
rect 83146 12218 83382 12454
rect 82826 11898 83062 12134
rect 83146 11898 83382 12134
rect 82826 -2502 83062 -2266
rect 83146 -2502 83382 -2266
rect 82826 -2822 83062 -2586
rect 83146 -2822 83382 -2586
rect 87326 707482 87562 707718
rect 87646 707482 87882 707718
rect 87326 707162 87562 707398
rect 87646 707162 87882 707398
rect 87326 700718 87562 700954
rect 87646 700718 87882 700954
rect 87326 700398 87562 700634
rect 87646 700398 87882 700634
rect 87326 664718 87562 664954
rect 87646 664718 87882 664954
rect 87326 664398 87562 664634
rect 87646 664398 87882 664634
rect 87326 628718 87562 628954
rect 87646 628718 87882 628954
rect 87326 628398 87562 628634
rect 87646 628398 87882 628634
rect 87326 592718 87562 592954
rect 87646 592718 87882 592954
rect 87326 592398 87562 592634
rect 87646 592398 87882 592634
rect 87326 556718 87562 556954
rect 87646 556718 87882 556954
rect 87326 556398 87562 556634
rect 87646 556398 87882 556634
rect 87326 520718 87562 520954
rect 87646 520718 87882 520954
rect 87326 520398 87562 520634
rect 87646 520398 87882 520634
rect 87326 484718 87562 484954
rect 87646 484718 87882 484954
rect 87326 484398 87562 484634
rect 87646 484398 87882 484634
rect 87326 448718 87562 448954
rect 87646 448718 87882 448954
rect 87326 448398 87562 448634
rect 87646 448398 87882 448634
rect 87326 412718 87562 412954
rect 87646 412718 87882 412954
rect 87326 412398 87562 412634
rect 87646 412398 87882 412634
rect 87326 376718 87562 376954
rect 87646 376718 87882 376954
rect 87326 376398 87562 376634
rect 87646 376398 87882 376634
rect 87326 340718 87562 340954
rect 87646 340718 87882 340954
rect 87326 340398 87562 340634
rect 87646 340398 87882 340634
rect 87326 304718 87562 304954
rect 87646 304718 87882 304954
rect 87326 304398 87562 304634
rect 87646 304398 87882 304634
rect 87326 268718 87562 268954
rect 87646 268718 87882 268954
rect 87326 268398 87562 268634
rect 87646 268398 87882 268634
rect 87326 232718 87562 232954
rect 87646 232718 87882 232954
rect 87326 232398 87562 232634
rect 87646 232398 87882 232634
rect 87326 196718 87562 196954
rect 87646 196718 87882 196954
rect 87326 196398 87562 196634
rect 87646 196398 87882 196634
rect 87326 160718 87562 160954
rect 87646 160718 87882 160954
rect 87326 160398 87562 160634
rect 87646 160398 87882 160634
rect 87326 124718 87562 124954
rect 87646 124718 87882 124954
rect 87326 124398 87562 124634
rect 87646 124398 87882 124634
rect 87326 88718 87562 88954
rect 87646 88718 87882 88954
rect 87326 88398 87562 88634
rect 87646 88398 87882 88634
rect 87326 52718 87562 52954
rect 87646 52718 87882 52954
rect 87326 52398 87562 52634
rect 87646 52398 87882 52634
rect 87326 16718 87562 16954
rect 87646 16718 87882 16954
rect 87326 16398 87562 16634
rect 87646 16398 87882 16634
rect 87326 -3462 87562 -3226
rect 87646 -3462 87882 -3226
rect 87326 -3782 87562 -3546
rect 87646 -3782 87882 -3546
rect 91826 708442 92062 708678
rect 92146 708442 92382 708678
rect 91826 708122 92062 708358
rect 92146 708122 92382 708358
rect 91826 669218 92062 669454
rect 92146 669218 92382 669454
rect 91826 668898 92062 669134
rect 92146 668898 92382 669134
rect 91826 633218 92062 633454
rect 92146 633218 92382 633454
rect 91826 632898 92062 633134
rect 92146 632898 92382 633134
rect 91826 597218 92062 597454
rect 92146 597218 92382 597454
rect 91826 596898 92062 597134
rect 92146 596898 92382 597134
rect 91826 561218 92062 561454
rect 92146 561218 92382 561454
rect 91826 560898 92062 561134
rect 92146 560898 92382 561134
rect 91826 525218 92062 525454
rect 92146 525218 92382 525454
rect 91826 524898 92062 525134
rect 92146 524898 92382 525134
rect 91826 489218 92062 489454
rect 92146 489218 92382 489454
rect 91826 488898 92062 489134
rect 92146 488898 92382 489134
rect 91826 453218 92062 453454
rect 92146 453218 92382 453454
rect 91826 452898 92062 453134
rect 92146 452898 92382 453134
rect 91826 417218 92062 417454
rect 92146 417218 92382 417454
rect 91826 416898 92062 417134
rect 92146 416898 92382 417134
rect 91826 381218 92062 381454
rect 92146 381218 92382 381454
rect 91826 380898 92062 381134
rect 92146 380898 92382 381134
rect 91826 345218 92062 345454
rect 92146 345218 92382 345454
rect 91826 344898 92062 345134
rect 92146 344898 92382 345134
rect 91826 309218 92062 309454
rect 92146 309218 92382 309454
rect 91826 308898 92062 309134
rect 92146 308898 92382 309134
rect 91826 273218 92062 273454
rect 92146 273218 92382 273454
rect 91826 272898 92062 273134
rect 92146 272898 92382 273134
rect 91826 237218 92062 237454
rect 92146 237218 92382 237454
rect 91826 236898 92062 237134
rect 92146 236898 92382 237134
rect 91826 201218 92062 201454
rect 92146 201218 92382 201454
rect 91826 200898 92062 201134
rect 92146 200898 92382 201134
rect 91826 165218 92062 165454
rect 92146 165218 92382 165454
rect 91826 164898 92062 165134
rect 92146 164898 92382 165134
rect 91826 129218 92062 129454
rect 92146 129218 92382 129454
rect 91826 128898 92062 129134
rect 92146 128898 92382 129134
rect 91826 93218 92062 93454
rect 92146 93218 92382 93454
rect 91826 92898 92062 93134
rect 92146 92898 92382 93134
rect 91826 57218 92062 57454
rect 92146 57218 92382 57454
rect 91826 56898 92062 57134
rect 92146 56898 92382 57134
rect 91826 21218 92062 21454
rect 92146 21218 92382 21454
rect 91826 20898 92062 21134
rect 92146 20898 92382 21134
rect 91826 -4422 92062 -4186
rect 92146 -4422 92382 -4186
rect 91826 -4742 92062 -4506
rect 92146 -4742 92382 -4506
rect 96326 709402 96562 709638
rect 96646 709402 96882 709638
rect 96326 709082 96562 709318
rect 96646 709082 96882 709318
rect 96326 673718 96562 673954
rect 96646 673718 96882 673954
rect 96326 673398 96562 673634
rect 96646 673398 96882 673634
rect 96326 637718 96562 637954
rect 96646 637718 96882 637954
rect 96326 637398 96562 637634
rect 96646 637398 96882 637634
rect 96326 601718 96562 601954
rect 96646 601718 96882 601954
rect 96326 601398 96562 601634
rect 96646 601398 96882 601634
rect 100826 710362 101062 710598
rect 101146 710362 101382 710598
rect 100826 710042 101062 710278
rect 101146 710042 101382 710278
rect 100826 678218 101062 678454
rect 101146 678218 101382 678454
rect 100826 677898 101062 678134
rect 101146 677898 101382 678134
rect 100826 642218 101062 642454
rect 101146 642218 101382 642454
rect 100826 641898 101062 642134
rect 101146 641898 101382 642134
rect 100826 606218 101062 606454
rect 101146 606218 101382 606454
rect 100826 605898 101062 606134
rect 101146 605898 101382 606134
rect 105326 711322 105562 711558
rect 105646 711322 105882 711558
rect 105326 711002 105562 711238
rect 105646 711002 105882 711238
rect 105326 682718 105562 682954
rect 105646 682718 105882 682954
rect 105326 682398 105562 682634
rect 105646 682398 105882 682634
rect 105326 646718 105562 646954
rect 105646 646718 105882 646954
rect 105326 646398 105562 646634
rect 105646 646398 105882 646634
rect 105326 610718 105562 610954
rect 105646 610718 105882 610954
rect 105326 610398 105562 610634
rect 105646 610398 105882 610634
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 109826 651218 110062 651454
rect 110146 651218 110382 651454
rect 109826 650898 110062 651134
rect 110146 650898 110382 651134
rect 109826 615218 110062 615454
rect 110146 615218 110382 615454
rect 109826 614898 110062 615134
rect 110146 614898 110382 615134
rect 114326 705562 114562 705798
rect 114646 705562 114882 705798
rect 114326 705242 114562 705478
rect 114646 705242 114882 705478
rect 114326 691718 114562 691954
rect 114646 691718 114882 691954
rect 114326 691398 114562 691634
rect 114646 691398 114882 691634
rect 114326 655718 114562 655954
rect 114646 655718 114882 655954
rect 114326 655398 114562 655634
rect 114646 655398 114882 655634
rect 114326 619718 114562 619954
rect 114646 619718 114882 619954
rect 114326 619398 114562 619634
rect 114646 619398 114882 619634
rect 118826 706522 119062 706758
rect 119146 706522 119382 706758
rect 118826 706202 119062 706438
rect 119146 706202 119382 706438
rect 118826 696218 119062 696454
rect 119146 696218 119382 696454
rect 118826 695898 119062 696134
rect 119146 695898 119382 696134
rect 118826 660218 119062 660454
rect 119146 660218 119382 660454
rect 118826 659898 119062 660134
rect 119146 659898 119382 660134
rect 118826 624218 119062 624454
rect 119146 624218 119382 624454
rect 118826 623898 119062 624134
rect 119146 623898 119382 624134
rect 123326 707482 123562 707718
rect 123646 707482 123882 707718
rect 123326 707162 123562 707398
rect 123646 707162 123882 707398
rect 123326 700718 123562 700954
rect 123646 700718 123882 700954
rect 123326 700398 123562 700634
rect 123646 700398 123882 700634
rect 123326 664718 123562 664954
rect 123646 664718 123882 664954
rect 123326 664398 123562 664634
rect 123646 664398 123882 664634
rect 123326 628718 123562 628954
rect 123646 628718 123882 628954
rect 123326 628398 123562 628634
rect 123646 628398 123882 628634
rect 123326 592718 123562 592954
rect 123646 592718 123882 592954
rect 123326 592398 123562 592634
rect 123646 592398 123882 592634
rect 127826 708442 128062 708678
rect 128146 708442 128382 708678
rect 127826 708122 128062 708358
rect 128146 708122 128382 708358
rect 127826 669218 128062 669454
rect 128146 669218 128382 669454
rect 127826 668898 128062 669134
rect 128146 668898 128382 669134
rect 127826 633218 128062 633454
rect 128146 633218 128382 633454
rect 127826 632898 128062 633134
rect 128146 632898 128382 633134
rect 127826 597218 128062 597454
rect 128146 597218 128382 597454
rect 127826 596898 128062 597134
rect 128146 596898 128382 597134
rect 132326 709402 132562 709638
rect 132646 709402 132882 709638
rect 132326 709082 132562 709318
rect 132646 709082 132882 709318
rect 132326 673718 132562 673954
rect 132646 673718 132882 673954
rect 132326 673398 132562 673634
rect 132646 673398 132882 673634
rect 132326 637718 132562 637954
rect 132646 637718 132882 637954
rect 132326 637398 132562 637634
rect 132646 637398 132882 637634
rect 132326 601718 132562 601954
rect 132646 601718 132882 601954
rect 132326 601398 132562 601634
rect 132646 601398 132882 601634
rect 136826 710362 137062 710598
rect 137146 710362 137382 710598
rect 136826 710042 137062 710278
rect 137146 710042 137382 710278
rect 136826 678218 137062 678454
rect 137146 678218 137382 678454
rect 136826 677898 137062 678134
rect 137146 677898 137382 678134
rect 136826 642218 137062 642454
rect 137146 642218 137382 642454
rect 136826 641898 137062 642134
rect 137146 641898 137382 642134
rect 136826 606218 137062 606454
rect 137146 606218 137382 606454
rect 136826 605898 137062 606134
rect 137146 605898 137382 606134
rect 141326 711322 141562 711558
rect 141646 711322 141882 711558
rect 141326 711002 141562 711238
rect 141646 711002 141882 711238
rect 141326 682718 141562 682954
rect 141646 682718 141882 682954
rect 141326 682398 141562 682634
rect 141646 682398 141882 682634
rect 141326 646718 141562 646954
rect 141646 646718 141882 646954
rect 141326 646398 141562 646634
rect 141646 646398 141882 646634
rect 141326 610718 141562 610954
rect 141646 610718 141882 610954
rect 141326 610398 141562 610634
rect 141646 610398 141882 610634
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 145826 651218 146062 651454
rect 146146 651218 146382 651454
rect 145826 650898 146062 651134
rect 146146 650898 146382 651134
rect 145826 615218 146062 615454
rect 146146 615218 146382 615454
rect 145826 614898 146062 615134
rect 146146 614898 146382 615134
rect 150326 705562 150562 705798
rect 150646 705562 150882 705798
rect 150326 705242 150562 705478
rect 150646 705242 150882 705478
rect 150326 691718 150562 691954
rect 150646 691718 150882 691954
rect 150326 691398 150562 691634
rect 150646 691398 150882 691634
rect 150326 655718 150562 655954
rect 150646 655718 150882 655954
rect 150326 655398 150562 655634
rect 150646 655398 150882 655634
rect 150326 619718 150562 619954
rect 150646 619718 150882 619954
rect 150326 619398 150562 619634
rect 150646 619398 150882 619634
rect 154826 706522 155062 706758
rect 155146 706522 155382 706758
rect 154826 706202 155062 706438
rect 155146 706202 155382 706438
rect 154826 696218 155062 696454
rect 155146 696218 155382 696454
rect 154826 695898 155062 696134
rect 155146 695898 155382 696134
rect 154826 660218 155062 660454
rect 155146 660218 155382 660454
rect 154826 659898 155062 660134
rect 155146 659898 155382 660134
rect 154826 624218 155062 624454
rect 155146 624218 155382 624454
rect 154826 623898 155062 624134
rect 155146 623898 155382 624134
rect 159326 707482 159562 707718
rect 159646 707482 159882 707718
rect 159326 707162 159562 707398
rect 159646 707162 159882 707398
rect 159326 700718 159562 700954
rect 159646 700718 159882 700954
rect 159326 700398 159562 700634
rect 159646 700398 159882 700634
rect 159326 664718 159562 664954
rect 159646 664718 159882 664954
rect 159326 664398 159562 664634
rect 159646 664398 159882 664634
rect 159326 628718 159562 628954
rect 159646 628718 159882 628954
rect 159326 628398 159562 628634
rect 159646 628398 159882 628634
rect 159326 592718 159562 592954
rect 159646 592718 159882 592954
rect 159326 592398 159562 592634
rect 159646 592398 159882 592634
rect 163826 708442 164062 708678
rect 164146 708442 164382 708678
rect 163826 708122 164062 708358
rect 164146 708122 164382 708358
rect 163826 669218 164062 669454
rect 164146 669218 164382 669454
rect 163826 668898 164062 669134
rect 164146 668898 164382 669134
rect 163826 633218 164062 633454
rect 164146 633218 164382 633454
rect 163826 632898 164062 633134
rect 164146 632898 164382 633134
rect 163826 597218 164062 597454
rect 164146 597218 164382 597454
rect 163826 596898 164062 597134
rect 164146 596898 164382 597134
rect 168326 709402 168562 709638
rect 168646 709402 168882 709638
rect 168326 709082 168562 709318
rect 168646 709082 168882 709318
rect 168326 673718 168562 673954
rect 168646 673718 168882 673954
rect 168326 673398 168562 673634
rect 168646 673398 168882 673634
rect 168326 637718 168562 637954
rect 168646 637718 168882 637954
rect 168326 637398 168562 637634
rect 168646 637398 168882 637634
rect 168326 601718 168562 601954
rect 168646 601718 168882 601954
rect 168326 601398 168562 601634
rect 168646 601398 168882 601634
rect 172826 710362 173062 710598
rect 173146 710362 173382 710598
rect 172826 710042 173062 710278
rect 173146 710042 173382 710278
rect 172826 678218 173062 678454
rect 173146 678218 173382 678454
rect 172826 677898 173062 678134
rect 173146 677898 173382 678134
rect 172826 642218 173062 642454
rect 173146 642218 173382 642454
rect 172826 641898 173062 642134
rect 173146 641898 173382 642134
rect 172826 606218 173062 606454
rect 173146 606218 173382 606454
rect 172826 605898 173062 606134
rect 173146 605898 173382 606134
rect 177326 711322 177562 711558
rect 177646 711322 177882 711558
rect 177326 711002 177562 711238
rect 177646 711002 177882 711238
rect 177326 682718 177562 682954
rect 177646 682718 177882 682954
rect 177326 682398 177562 682634
rect 177646 682398 177882 682634
rect 177326 646718 177562 646954
rect 177646 646718 177882 646954
rect 177326 646398 177562 646634
rect 177646 646398 177882 646634
rect 177326 610718 177562 610954
rect 177646 610718 177882 610954
rect 177326 610398 177562 610634
rect 177646 610398 177882 610634
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 181826 651218 182062 651454
rect 182146 651218 182382 651454
rect 181826 650898 182062 651134
rect 182146 650898 182382 651134
rect 181826 615218 182062 615454
rect 182146 615218 182382 615454
rect 181826 614898 182062 615134
rect 182146 614898 182382 615134
rect 186326 705562 186562 705798
rect 186646 705562 186882 705798
rect 186326 705242 186562 705478
rect 186646 705242 186882 705478
rect 186326 691718 186562 691954
rect 186646 691718 186882 691954
rect 186326 691398 186562 691634
rect 186646 691398 186882 691634
rect 186326 655718 186562 655954
rect 186646 655718 186882 655954
rect 186326 655398 186562 655634
rect 186646 655398 186882 655634
rect 186326 619718 186562 619954
rect 186646 619718 186882 619954
rect 186326 619398 186562 619634
rect 186646 619398 186882 619634
rect 190826 706522 191062 706758
rect 191146 706522 191382 706758
rect 190826 706202 191062 706438
rect 191146 706202 191382 706438
rect 190826 696218 191062 696454
rect 191146 696218 191382 696454
rect 190826 695898 191062 696134
rect 191146 695898 191382 696134
rect 190826 660218 191062 660454
rect 191146 660218 191382 660454
rect 190826 659898 191062 660134
rect 191146 659898 191382 660134
rect 190826 624218 191062 624454
rect 191146 624218 191382 624454
rect 190826 623898 191062 624134
rect 191146 623898 191382 624134
rect 195326 707482 195562 707718
rect 195646 707482 195882 707718
rect 195326 707162 195562 707398
rect 195646 707162 195882 707398
rect 195326 700718 195562 700954
rect 195646 700718 195882 700954
rect 195326 700398 195562 700634
rect 195646 700398 195882 700634
rect 195326 664718 195562 664954
rect 195646 664718 195882 664954
rect 195326 664398 195562 664634
rect 195646 664398 195882 664634
rect 195326 628718 195562 628954
rect 195646 628718 195882 628954
rect 195326 628398 195562 628634
rect 195646 628398 195882 628634
rect 195326 592718 195562 592954
rect 195646 592718 195882 592954
rect 195326 592398 195562 592634
rect 195646 592398 195882 592634
rect 100328 583718 100564 583954
rect 100328 583398 100564 583634
rect 190496 583718 190732 583954
rect 190496 583398 190732 583634
rect 101008 579218 101244 579454
rect 101008 578898 101244 579134
rect 189816 579218 190052 579454
rect 189816 578898 190052 579134
rect 96326 565718 96562 565954
rect 96646 565718 96882 565954
rect 96326 565398 96562 565634
rect 96646 565398 96882 565634
rect 195326 556718 195562 556954
rect 195646 556718 195882 556954
rect 195326 556398 195562 556634
rect 195646 556398 195882 556634
rect 100328 547718 100564 547954
rect 100328 547398 100564 547634
rect 190496 547718 190732 547954
rect 190496 547398 190732 547634
rect 101008 543218 101244 543454
rect 101008 542898 101244 543134
rect 189816 543218 190052 543454
rect 189816 542898 190052 543134
rect 96326 529718 96562 529954
rect 96646 529718 96882 529954
rect 96326 529398 96562 529634
rect 96646 529398 96882 529634
rect 195326 520718 195562 520954
rect 195646 520718 195882 520954
rect 195326 520398 195562 520634
rect 195646 520398 195882 520634
rect 100328 511718 100564 511954
rect 100328 511398 100564 511634
rect 190496 511718 190732 511954
rect 190496 511398 190732 511634
rect 101008 507218 101244 507454
rect 101008 506898 101244 507134
rect 189816 507218 190052 507454
rect 189816 506898 190052 507134
rect 96326 493718 96562 493954
rect 96646 493718 96882 493954
rect 96326 493398 96562 493634
rect 96646 493398 96882 493634
rect 96326 457718 96562 457954
rect 96646 457718 96882 457954
rect 96326 457398 96562 457634
rect 96646 457398 96882 457634
rect 96326 421718 96562 421954
rect 96646 421718 96882 421954
rect 96326 421398 96562 421634
rect 96646 421398 96882 421634
rect 96326 385718 96562 385954
rect 96646 385718 96882 385954
rect 96326 385398 96562 385634
rect 96646 385398 96882 385634
rect 96326 349718 96562 349954
rect 96646 349718 96882 349954
rect 96326 349398 96562 349634
rect 96646 349398 96882 349634
rect 96326 313718 96562 313954
rect 96646 313718 96882 313954
rect 96326 313398 96562 313634
rect 96646 313398 96882 313634
rect 96326 277718 96562 277954
rect 96646 277718 96882 277954
rect 96326 277398 96562 277634
rect 96646 277398 96882 277634
rect 96326 241718 96562 241954
rect 96646 241718 96882 241954
rect 96326 241398 96562 241634
rect 96646 241398 96882 241634
rect 96326 205718 96562 205954
rect 96646 205718 96882 205954
rect 96326 205398 96562 205634
rect 96646 205398 96882 205634
rect 96326 169718 96562 169954
rect 96646 169718 96882 169954
rect 96326 169398 96562 169634
rect 96646 169398 96882 169634
rect 96326 133718 96562 133954
rect 96646 133718 96882 133954
rect 96326 133398 96562 133634
rect 96646 133398 96882 133634
rect 96326 97718 96562 97954
rect 96646 97718 96882 97954
rect 96326 97398 96562 97634
rect 96646 97398 96882 97634
rect 96326 61718 96562 61954
rect 96646 61718 96882 61954
rect 96326 61398 96562 61634
rect 96646 61398 96882 61634
rect 96326 25718 96562 25954
rect 96646 25718 96882 25954
rect 96326 25398 96562 25634
rect 96646 25398 96882 25634
rect 96326 -5382 96562 -5146
rect 96646 -5382 96882 -5146
rect 96326 -5702 96562 -5466
rect 96646 -5702 96882 -5466
rect 100826 462218 101062 462454
rect 101146 462218 101382 462454
rect 100826 461898 101062 462134
rect 101146 461898 101382 462134
rect 100826 426218 101062 426454
rect 101146 426218 101382 426454
rect 100826 425898 101062 426134
rect 101146 425898 101382 426134
rect 100826 390218 101062 390454
rect 101146 390218 101382 390454
rect 100826 389898 101062 390134
rect 101146 389898 101382 390134
rect 100826 354218 101062 354454
rect 101146 354218 101382 354454
rect 100826 353898 101062 354134
rect 101146 353898 101382 354134
rect 100826 318218 101062 318454
rect 101146 318218 101382 318454
rect 100826 317898 101062 318134
rect 101146 317898 101382 318134
rect 100826 282218 101062 282454
rect 101146 282218 101382 282454
rect 100826 281898 101062 282134
rect 101146 281898 101382 282134
rect 100826 246218 101062 246454
rect 101146 246218 101382 246454
rect 100826 245898 101062 246134
rect 101146 245898 101382 246134
rect 100826 210218 101062 210454
rect 101146 210218 101382 210454
rect 100826 209898 101062 210134
rect 101146 209898 101382 210134
rect 100826 174218 101062 174454
rect 101146 174218 101382 174454
rect 100826 173898 101062 174134
rect 101146 173898 101382 174134
rect 100826 138218 101062 138454
rect 101146 138218 101382 138454
rect 100826 137898 101062 138134
rect 101146 137898 101382 138134
rect 100826 102218 101062 102454
rect 101146 102218 101382 102454
rect 100826 101898 101062 102134
rect 101146 101898 101382 102134
rect 100826 66218 101062 66454
rect 101146 66218 101382 66454
rect 100826 65898 101062 66134
rect 101146 65898 101382 66134
rect 100826 30218 101062 30454
rect 101146 30218 101382 30454
rect 100826 29898 101062 30134
rect 101146 29898 101382 30134
rect 100826 -6342 101062 -6106
rect 101146 -6342 101382 -6106
rect 100826 -6662 101062 -6426
rect 101146 -6662 101382 -6426
rect 105326 466718 105562 466954
rect 105646 466718 105882 466954
rect 105326 466398 105562 466634
rect 105646 466398 105882 466634
rect 105326 430718 105562 430954
rect 105646 430718 105882 430954
rect 105326 430398 105562 430634
rect 105646 430398 105882 430634
rect 105326 394718 105562 394954
rect 105646 394718 105882 394954
rect 105326 394398 105562 394634
rect 105646 394398 105882 394634
rect 105326 358718 105562 358954
rect 105646 358718 105882 358954
rect 105326 358398 105562 358634
rect 105646 358398 105882 358634
rect 105326 322718 105562 322954
rect 105646 322718 105882 322954
rect 105326 322398 105562 322634
rect 105646 322398 105882 322634
rect 105326 286718 105562 286954
rect 105646 286718 105882 286954
rect 105326 286398 105562 286634
rect 105646 286398 105882 286634
rect 105326 250718 105562 250954
rect 105646 250718 105882 250954
rect 105326 250398 105562 250634
rect 105646 250398 105882 250634
rect 105326 214718 105562 214954
rect 105646 214718 105882 214954
rect 105326 214398 105562 214634
rect 105646 214398 105882 214634
rect 105326 178718 105562 178954
rect 105646 178718 105882 178954
rect 105326 178398 105562 178634
rect 105646 178398 105882 178634
rect 105326 142718 105562 142954
rect 105646 142718 105882 142954
rect 105326 142398 105562 142634
rect 105646 142398 105882 142634
rect 105326 106718 105562 106954
rect 105646 106718 105882 106954
rect 105326 106398 105562 106634
rect 105646 106398 105882 106634
rect 105326 70718 105562 70954
rect 105646 70718 105882 70954
rect 105326 70398 105562 70634
rect 105646 70398 105882 70634
rect 105326 34718 105562 34954
rect 105646 34718 105882 34954
rect 105326 34398 105562 34634
rect 105646 34398 105882 34634
rect 105326 -7302 105562 -7066
rect 105646 -7302 105882 -7066
rect 105326 -7622 105562 -7386
rect 105646 -7622 105882 -7386
rect 109826 471218 110062 471454
rect 110146 471218 110382 471454
rect 109826 470898 110062 471134
rect 110146 470898 110382 471134
rect 109826 435218 110062 435454
rect 110146 435218 110382 435454
rect 109826 434898 110062 435134
rect 110146 434898 110382 435134
rect 109826 399218 110062 399454
rect 110146 399218 110382 399454
rect 109826 398898 110062 399134
rect 110146 398898 110382 399134
rect 109826 363218 110062 363454
rect 110146 363218 110382 363454
rect 109826 362898 110062 363134
rect 110146 362898 110382 363134
rect 109826 327218 110062 327454
rect 110146 327218 110382 327454
rect 109826 326898 110062 327134
rect 110146 326898 110382 327134
rect 109826 291218 110062 291454
rect 110146 291218 110382 291454
rect 109826 290898 110062 291134
rect 110146 290898 110382 291134
rect 109826 255218 110062 255454
rect 110146 255218 110382 255454
rect 109826 254898 110062 255134
rect 110146 254898 110382 255134
rect 109826 219218 110062 219454
rect 110146 219218 110382 219454
rect 109826 218898 110062 219134
rect 110146 218898 110382 219134
rect 109826 183218 110062 183454
rect 110146 183218 110382 183454
rect 109826 182898 110062 183134
rect 110146 182898 110382 183134
rect 109826 147218 110062 147454
rect 110146 147218 110382 147454
rect 109826 146898 110062 147134
rect 110146 146898 110382 147134
rect 109826 111218 110062 111454
rect 110146 111218 110382 111454
rect 109826 110898 110062 111134
rect 110146 110898 110382 111134
rect 109826 75218 110062 75454
rect 110146 75218 110382 75454
rect 109826 74898 110062 75134
rect 110146 74898 110382 75134
rect 109826 39218 110062 39454
rect 110146 39218 110382 39454
rect 109826 38898 110062 39134
rect 110146 38898 110382 39134
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 114326 475718 114562 475954
rect 114646 475718 114882 475954
rect 114326 475398 114562 475634
rect 114646 475398 114882 475634
rect 114326 439718 114562 439954
rect 114646 439718 114882 439954
rect 114326 439398 114562 439634
rect 114646 439398 114882 439634
rect 114326 403718 114562 403954
rect 114646 403718 114882 403954
rect 114326 403398 114562 403634
rect 114646 403398 114882 403634
rect 114326 367718 114562 367954
rect 114646 367718 114882 367954
rect 114326 367398 114562 367634
rect 114646 367398 114882 367634
rect 114326 331718 114562 331954
rect 114646 331718 114882 331954
rect 114326 331398 114562 331634
rect 114646 331398 114882 331634
rect 114326 295718 114562 295954
rect 114646 295718 114882 295954
rect 114326 295398 114562 295634
rect 114646 295398 114882 295634
rect 114326 259718 114562 259954
rect 114646 259718 114882 259954
rect 114326 259398 114562 259634
rect 114646 259398 114882 259634
rect 114326 223718 114562 223954
rect 114646 223718 114882 223954
rect 114326 223398 114562 223634
rect 114646 223398 114882 223634
rect 114326 187718 114562 187954
rect 114646 187718 114882 187954
rect 114326 187398 114562 187634
rect 114646 187398 114882 187634
rect 114326 151718 114562 151954
rect 114646 151718 114882 151954
rect 114326 151398 114562 151634
rect 114646 151398 114882 151634
rect 114326 115718 114562 115954
rect 114646 115718 114882 115954
rect 114326 115398 114562 115634
rect 114646 115398 114882 115634
rect 114326 79718 114562 79954
rect 114646 79718 114882 79954
rect 114326 79398 114562 79634
rect 114646 79398 114882 79634
rect 114326 43718 114562 43954
rect 114646 43718 114882 43954
rect 114326 43398 114562 43634
rect 114646 43398 114882 43634
rect 114326 7718 114562 7954
rect 114646 7718 114882 7954
rect 114326 7398 114562 7634
rect 114646 7398 114882 7634
rect 114326 -1542 114562 -1306
rect 114646 -1542 114882 -1306
rect 114326 -1862 114562 -1626
rect 114646 -1862 114882 -1626
rect 118826 480218 119062 480454
rect 119146 480218 119382 480454
rect 118826 479898 119062 480134
rect 119146 479898 119382 480134
rect 118826 444218 119062 444454
rect 119146 444218 119382 444454
rect 118826 443898 119062 444134
rect 119146 443898 119382 444134
rect 118826 408218 119062 408454
rect 119146 408218 119382 408454
rect 118826 407898 119062 408134
rect 119146 407898 119382 408134
rect 118826 372218 119062 372454
rect 119146 372218 119382 372454
rect 118826 371898 119062 372134
rect 119146 371898 119382 372134
rect 118826 336218 119062 336454
rect 119146 336218 119382 336454
rect 118826 335898 119062 336134
rect 119146 335898 119382 336134
rect 118826 300218 119062 300454
rect 119146 300218 119382 300454
rect 118826 299898 119062 300134
rect 119146 299898 119382 300134
rect 118826 264218 119062 264454
rect 119146 264218 119382 264454
rect 118826 263898 119062 264134
rect 119146 263898 119382 264134
rect 118826 228218 119062 228454
rect 119146 228218 119382 228454
rect 118826 227898 119062 228134
rect 119146 227898 119382 228134
rect 118826 192218 119062 192454
rect 119146 192218 119382 192454
rect 118826 191898 119062 192134
rect 119146 191898 119382 192134
rect 118826 156218 119062 156454
rect 119146 156218 119382 156454
rect 118826 155898 119062 156134
rect 119146 155898 119382 156134
rect 118826 120218 119062 120454
rect 119146 120218 119382 120454
rect 118826 119898 119062 120134
rect 119146 119898 119382 120134
rect 118826 84218 119062 84454
rect 119146 84218 119382 84454
rect 118826 83898 119062 84134
rect 119146 83898 119382 84134
rect 118826 48218 119062 48454
rect 119146 48218 119382 48454
rect 118826 47898 119062 48134
rect 119146 47898 119382 48134
rect 118826 12218 119062 12454
rect 119146 12218 119382 12454
rect 118826 11898 119062 12134
rect 119146 11898 119382 12134
rect 118826 -2502 119062 -2266
rect 119146 -2502 119382 -2266
rect 118826 -2822 119062 -2586
rect 119146 -2822 119382 -2586
rect 123326 484718 123562 484954
rect 123646 484718 123882 484954
rect 123326 484398 123562 484634
rect 123646 484398 123882 484634
rect 123326 448718 123562 448954
rect 123646 448718 123882 448954
rect 123326 448398 123562 448634
rect 123646 448398 123882 448634
rect 123326 412718 123562 412954
rect 123646 412718 123882 412954
rect 123326 412398 123562 412634
rect 123646 412398 123882 412634
rect 123326 376718 123562 376954
rect 123646 376718 123882 376954
rect 123326 376398 123562 376634
rect 123646 376398 123882 376634
rect 123326 340718 123562 340954
rect 123646 340718 123882 340954
rect 123326 340398 123562 340634
rect 123646 340398 123882 340634
rect 123326 304718 123562 304954
rect 123646 304718 123882 304954
rect 123326 304398 123562 304634
rect 123646 304398 123882 304634
rect 123326 268718 123562 268954
rect 123646 268718 123882 268954
rect 123326 268398 123562 268634
rect 123646 268398 123882 268634
rect 123326 232718 123562 232954
rect 123646 232718 123882 232954
rect 123326 232398 123562 232634
rect 123646 232398 123882 232634
rect 123326 196718 123562 196954
rect 123646 196718 123882 196954
rect 123326 196398 123562 196634
rect 123646 196398 123882 196634
rect 123326 160718 123562 160954
rect 123646 160718 123882 160954
rect 123326 160398 123562 160634
rect 123646 160398 123882 160634
rect 123326 124718 123562 124954
rect 123646 124718 123882 124954
rect 123326 124398 123562 124634
rect 123646 124398 123882 124634
rect 123326 88718 123562 88954
rect 123646 88718 123882 88954
rect 123326 88398 123562 88634
rect 123646 88398 123882 88634
rect 123326 52718 123562 52954
rect 123646 52718 123882 52954
rect 123326 52398 123562 52634
rect 123646 52398 123882 52634
rect 123326 16718 123562 16954
rect 123646 16718 123882 16954
rect 123326 16398 123562 16634
rect 123646 16398 123882 16634
rect 123326 -3462 123562 -3226
rect 123646 -3462 123882 -3226
rect 123326 -3782 123562 -3546
rect 123646 -3782 123882 -3546
rect 127826 489218 128062 489454
rect 128146 489218 128382 489454
rect 127826 488898 128062 489134
rect 128146 488898 128382 489134
rect 127826 453218 128062 453454
rect 128146 453218 128382 453454
rect 127826 452898 128062 453134
rect 128146 452898 128382 453134
rect 127826 417218 128062 417454
rect 128146 417218 128382 417454
rect 127826 416898 128062 417134
rect 128146 416898 128382 417134
rect 127826 381218 128062 381454
rect 128146 381218 128382 381454
rect 127826 380898 128062 381134
rect 128146 380898 128382 381134
rect 127826 345218 128062 345454
rect 128146 345218 128382 345454
rect 127826 344898 128062 345134
rect 128146 344898 128382 345134
rect 127826 309218 128062 309454
rect 128146 309218 128382 309454
rect 127826 308898 128062 309134
rect 128146 308898 128382 309134
rect 127826 273218 128062 273454
rect 128146 273218 128382 273454
rect 127826 272898 128062 273134
rect 128146 272898 128382 273134
rect 127826 237218 128062 237454
rect 128146 237218 128382 237454
rect 127826 236898 128062 237134
rect 128146 236898 128382 237134
rect 127826 201218 128062 201454
rect 128146 201218 128382 201454
rect 127826 200898 128062 201134
rect 128146 200898 128382 201134
rect 127826 165218 128062 165454
rect 128146 165218 128382 165454
rect 127826 164898 128062 165134
rect 128146 164898 128382 165134
rect 127826 129218 128062 129454
rect 128146 129218 128382 129454
rect 127826 128898 128062 129134
rect 128146 128898 128382 129134
rect 127826 93218 128062 93454
rect 128146 93218 128382 93454
rect 127826 92898 128062 93134
rect 128146 92898 128382 93134
rect 127826 57218 128062 57454
rect 128146 57218 128382 57454
rect 127826 56898 128062 57134
rect 128146 56898 128382 57134
rect 127826 21218 128062 21454
rect 128146 21218 128382 21454
rect 127826 20898 128062 21134
rect 128146 20898 128382 21134
rect 127826 -4422 128062 -4186
rect 128146 -4422 128382 -4186
rect 127826 -4742 128062 -4506
rect 128146 -4742 128382 -4506
rect 132326 493718 132562 493954
rect 132646 493718 132882 493954
rect 132326 493398 132562 493634
rect 132646 493398 132882 493634
rect 132326 457718 132562 457954
rect 132646 457718 132882 457954
rect 132326 457398 132562 457634
rect 132646 457398 132882 457634
rect 132326 421718 132562 421954
rect 132646 421718 132882 421954
rect 132326 421398 132562 421634
rect 132646 421398 132882 421634
rect 132326 385718 132562 385954
rect 132646 385718 132882 385954
rect 132326 385398 132562 385634
rect 132646 385398 132882 385634
rect 132326 349718 132562 349954
rect 132646 349718 132882 349954
rect 132326 349398 132562 349634
rect 132646 349398 132882 349634
rect 132326 313718 132562 313954
rect 132646 313718 132882 313954
rect 132326 313398 132562 313634
rect 132646 313398 132882 313634
rect 132326 277718 132562 277954
rect 132646 277718 132882 277954
rect 132326 277398 132562 277634
rect 132646 277398 132882 277634
rect 132326 241718 132562 241954
rect 132646 241718 132882 241954
rect 132326 241398 132562 241634
rect 132646 241398 132882 241634
rect 132326 205718 132562 205954
rect 132646 205718 132882 205954
rect 132326 205398 132562 205634
rect 132646 205398 132882 205634
rect 132326 169718 132562 169954
rect 132646 169718 132882 169954
rect 132326 169398 132562 169634
rect 132646 169398 132882 169634
rect 132326 133718 132562 133954
rect 132646 133718 132882 133954
rect 132326 133398 132562 133634
rect 132646 133398 132882 133634
rect 132326 97718 132562 97954
rect 132646 97718 132882 97954
rect 132326 97398 132562 97634
rect 132646 97398 132882 97634
rect 132326 61718 132562 61954
rect 132646 61718 132882 61954
rect 132326 61398 132562 61634
rect 132646 61398 132882 61634
rect 132326 25718 132562 25954
rect 132646 25718 132882 25954
rect 132326 25398 132562 25634
rect 132646 25398 132882 25634
rect 132326 -5382 132562 -5146
rect 132646 -5382 132882 -5146
rect 132326 -5702 132562 -5466
rect 132646 -5702 132882 -5466
rect 136826 462218 137062 462454
rect 137146 462218 137382 462454
rect 136826 461898 137062 462134
rect 137146 461898 137382 462134
rect 136826 426218 137062 426454
rect 137146 426218 137382 426454
rect 136826 425898 137062 426134
rect 137146 425898 137382 426134
rect 136826 390218 137062 390454
rect 137146 390218 137382 390454
rect 136826 389898 137062 390134
rect 137146 389898 137382 390134
rect 136826 354218 137062 354454
rect 137146 354218 137382 354454
rect 136826 353898 137062 354134
rect 137146 353898 137382 354134
rect 136826 318218 137062 318454
rect 137146 318218 137382 318454
rect 136826 317898 137062 318134
rect 137146 317898 137382 318134
rect 136826 282218 137062 282454
rect 137146 282218 137382 282454
rect 136826 281898 137062 282134
rect 137146 281898 137382 282134
rect 136826 246218 137062 246454
rect 137146 246218 137382 246454
rect 136826 245898 137062 246134
rect 137146 245898 137382 246134
rect 136826 210218 137062 210454
rect 137146 210218 137382 210454
rect 136826 209898 137062 210134
rect 137146 209898 137382 210134
rect 136826 174218 137062 174454
rect 137146 174218 137382 174454
rect 136826 173898 137062 174134
rect 137146 173898 137382 174134
rect 136826 138218 137062 138454
rect 137146 138218 137382 138454
rect 136826 137898 137062 138134
rect 137146 137898 137382 138134
rect 136826 102218 137062 102454
rect 137146 102218 137382 102454
rect 136826 101898 137062 102134
rect 137146 101898 137382 102134
rect 136826 66218 137062 66454
rect 137146 66218 137382 66454
rect 136826 65898 137062 66134
rect 137146 65898 137382 66134
rect 136826 30218 137062 30454
rect 137146 30218 137382 30454
rect 136826 29898 137062 30134
rect 137146 29898 137382 30134
rect 136826 -6342 137062 -6106
rect 137146 -6342 137382 -6106
rect 136826 -6662 137062 -6426
rect 137146 -6662 137382 -6426
rect 141326 466718 141562 466954
rect 141646 466718 141882 466954
rect 141326 466398 141562 466634
rect 141646 466398 141882 466634
rect 141326 430718 141562 430954
rect 141646 430718 141882 430954
rect 141326 430398 141562 430634
rect 141646 430398 141882 430634
rect 141326 394718 141562 394954
rect 141646 394718 141882 394954
rect 141326 394398 141562 394634
rect 141646 394398 141882 394634
rect 141326 358718 141562 358954
rect 141646 358718 141882 358954
rect 141326 358398 141562 358634
rect 141646 358398 141882 358634
rect 141326 322718 141562 322954
rect 141646 322718 141882 322954
rect 141326 322398 141562 322634
rect 141646 322398 141882 322634
rect 141326 286718 141562 286954
rect 141646 286718 141882 286954
rect 141326 286398 141562 286634
rect 141646 286398 141882 286634
rect 141326 250718 141562 250954
rect 141646 250718 141882 250954
rect 141326 250398 141562 250634
rect 141646 250398 141882 250634
rect 141326 214718 141562 214954
rect 141646 214718 141882 214954
rect 141326 214398 141562 214634
rect 141646 214398 141882 214634
rect 141326 178718 141562 178954
rect 141646 178718 141882 178954
rect 141326 178398 141562 178634
rect 141646 178398 141882 178634
rect 141326 142718 141562 142954
rect 141646 142718 141882 142954
rect 141326 142398 141562 142634
rect 141646 142398 141882 142634
rect 141326 106718 141562 106954
rect 141646 106718 141882 106954
rect 141326 106398 141562 106634
rect 141646 106398 141882 106634
rect 141326 70718 141562 70954
rect 141646 70718 141882 70954
rect 141326 70398 141562 70634
rect 141646 70398 141882 70634
rect 141326 34718 141562 34954
rect 141646 34718 141882 34954
rect 141326 34398 141562 34634
rect 141646 34398 141882 34634
rect 141326 -7302 141562 -7066
rect 141646 -7302 141882 -7066
rect 141326 -7622 141562 -7386
rect 141646 -7622 141882 -7386
rect 145826 471218 146062 471454
rect 146146 471218 146382 471454
rect 145826 470898 146062 471134
rect 146146 470898 146382 471134
rect 145826 435218 146062 435454
rect 146146 435218 146382 435454
rect 145826 434898 146062 435134
rect 146146 434898 146382 435134
rect 145826 399218 146062 399454
rect 146146 399218 146382 399454
rect 145826 398898 146062 399134
rect 146146 398898 146382 399134
rect 145826 363218 146062 363454
rect 146146 363218 146382 363454
rect 145826 362898 146062 363134
rect 146146 362898 146382 363134
rect 145826 327218 146062 327454
rect 146146 327218 146382 327454
rect 145826 326898 146062 327134
rect 146146 326898 146382 327134
rect 145826 291218 146062 291454
rect 146146 291218 146382 291454
rect 145826 290898 146062 291134
rect 146146 290898 146382 291134
rect 145826 255218 146062 255454
rect 146146 255218 146382 255454
rect 145826 254898 146062 255134
rect 146146 254898 146382 255134
rect 145826 219218 146062 219454
rect 146146 219218 146382 219454
rect 145826 218898 146062 219134
rect 146146 218898 146382 219134
rect 145826 183218 146062 183454
rect 146146 183218 146382 183454
rect 145826 182898 146062 183134
rect 146146 182898 146382 183134
rect 145826 147218 146062 147454
rect 146146 147218 146382 147454
rect 145826 146898 146062 147134
rect 146146 146898 146382 147134
rect 145826 111218 146062 111454
rect 146146 111218 146382 111454
rect 145826 110898 146062 111134
rect 146146 110898 146382 111134
rect 145826 75218 146062 75454
rect 146146 75218 146382 75454
rect 145826 74898 146062 75134
rect 146146 74898 146382 75134
rect 145826 39218 146062 39454
rect 146146 39218 146382 39454
rect 145826 38898 146062 39134
rect 146146 38898 146382 39134
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 150326 475718 150562 475954
rect 150646 475718 150882 475954
rect 150326 475398 150562 475634
rect 150646 475398 150882 475634
rect 150326 439718 150562 439954
rect 150646 439718 150882 439954
rect 150326 439398 150562 439634
rect 150646 439398 150882 439634
rect 150326 403718 150562 403954
rect 150646 403718 150882 403954
rect 150326 403398 150562 403634
rect 150646 403398 150882 403634
rect 150326 367718 150562 367954
rect 150646 367718 150882 367954
rect 150326 367398 150562 367634
rect 150646 367398 150882 367634
rect 150326 331718 150562 331954
rect 150646 331718 150882 331954
rect 150326 331398 150562 331634
rect 150646 331398 150882 331634
rect 150326 295718 150562 295954
rect 150646 295718 150882 295954
rect 150326 295398 150562 295634
rect 150646 295398 150882 295634
rect 150326 259718 150562 259954
rect 150646 259718 150882 259954
rect 150326 259398 150562 259634
rect 150646 259398 150882 259634
rect 150326 223718 150562 223954
rect 150646 223718 150882 223954
rect 150326 223398 150562 223634
rect 150646 223398 150882 223634
rect 150326 187718 150562 187954
rect 150646 187718 150882 187954
rect 150326 187398 150562 187634
rect 150646 187398 150882 187634
rect 150326 151718 150562 151954
rect 150646 151718 150882 151954
rect 150326 151398 150562 151634
rect 150646 151398 150882 151634
rect 150326 115718 150562 115954
rect 150646 115718 150882 115954
rect 150326 115398 150562 115634
rect 150646 115398 150882 115634
rect 150326 79718 150562 79954
rect 150646 79718 150882 79954
rect 150326 79398 150562 79634
rect 150646 79398 150882 79634
rect 150326 43718 150562 43954
rect 150646 43718 150882 43954
rect 150326 43398 150562 43634
rect 150646 43398 150882 43634
rect 150326 7718 150562 7954
rect 150646 7718 150882 7954
rect 150326 7398 150562 7634
rect 150646 7398 150882 7634
rect 150326 -1542 150562 -1306
rect 150646 -1542 150882 -1306
rect 150326 -1862 150562 -1626
rect 150646 -1862 150882 -1626
rect 154826 480218 155062 480454
rect 155146 480218 155382 480454
rect 154826 479898 155062 480134
rect 155146 479898 155382 480134
rect 154826 444218 155062 444454
rect 155146 444218 155382 444454
rect 154826 443898 155062 444134
rect 155146 443898 155382 444134
rect 154826 408218 155062 408454
rect 155146 408218 155382 408454
rect 154826 407898 155062 408134
rect 155146 407898 155382 408134
rect 154826 372218 155062 372454
rect 155146 372218 155382 372454
rect 154826 371898 155062 372134
rect 155146 371898 155382 372134
rect 154826 336218 155062 336454
rect 155146 336218 155382 336454
rect 154826 335898 155062 336134
rect 155146 335898 155382 336134
rect 154826 300218 155062 300454
rect 155146 300218 155382 300454
rect 154826 299898 155062 300134
rect 155146 299898 155382 300134
rect 154826 264218 155062 264454
rect 155146 264218 155382 264454
rect 154826 263898 155062 264134
rect 155146 263898 155382 264134
rect 154826 228218 155062 228454
rect 155146 228218 155382 228454
rect 154826 227898 155062 228134
rect 155146 227898 155382 228134
rect 154826 192218 155062 192454
rect 155146 192218 155382 192454
rect 154826 191898 155062 192134
rect 155146 191898 155382 192134
rect 154826 156218 155062 156454
rect 155146 156218 155382 156454
rect 154826 155898 155062 156134
rect 155146 155898 155382 156134
rect 154826 120218 155062 120454
rect 155146 120218 155382 120454
rect 154826 119898 155062 120134
rect 155146 119898 155382 120134
rect 154826 84218 155062 84454
rect 155146 84218 155382 84454
rect 154826 83898 155062 84134
rect 155146 83898 155382 84134
rect 154826 48218 155062 48454
rect 155146 48218 155382 48454
rect 154826 47898 155062 48134
rect 155146 47898 155382 48134
rect 154826 12218 155062 12454
rect 155146 12218 155382 12454
rect 154826 11898 155062 12134
rect 155146 11898 155382 12134
rect 154826 -2502 155062 -2266
rect 155146 -2502 155382 -2266
rect 154826 -2822 155062 -2586
rect 155146 -2822 155382 -2586
rect 159326 484718 159562 484954
rect 159646 484718 159882 484954
rect 159326 484398 159562 484634
rect 159646 484398 159882 484634
rect 159326 448718 159562 448954
rect 159646 448718 159882 448954
rect 159326 448398 159562 448634
rect 159646 448398 159882 448634
rect 159326 412718 159562 412954
rect 159646 412718 159882 412954
rect 159326 412398 159562 412634
rect 159646 412398 159882 412634
rect 159326 376718 159562 376954
rect 159646 376718 159882 376954
rect 159326 376398 159562 376634
rect 159646 376398 159882 376634
rect 159326 340718 159562 340954
rect 159646 340718 159882 340954
rect 159326 340398 159562 340634
rect 159646 340398 159882 340634
rect 159326 304718 159562 304954
rect 159646 304718 159882 304954
rect 159326 304398 159562 304634
rect 159646 304398 159882 304634
rect 159326 268718 159562 268954
rect 159646 268718 159882 268954
rect 159326 268398 159562 268634
rect 159646 268398 159882 268634
rect 159326 232718 159562 232954
rect 159646 232718 159882 232954
rect 159326 232398 159562 232634
rect 159646 232398 159882 232634
rect 159326 196718 159562 196954
rect 159646 196718 159882 196954
rect 159326 196398 159562 196634
rect 159646 196398 159882 196634
rect 159326 160718 159562 160954
rect 159646 160718 159882 160954
rect 159326 160398 159562 160634
rect 159646 160398 159882 160634
rect 159326 124718 159562 124954
rect 159646 124718 159882 124954
rect 159326 124398 159562 124634
rect 159646 124398 159882 124634
rect 159326 88718 159562 88954
rect 159646 88718 159882 88954
rect 159326 88398 159562 88634
rect 159646 88398 159882 88634
rect 159326 52718 159562 52954
rect 159646 52718 159882 52954
rect 159326 52398 159562 52634
rect 159646 52398 159882 52634
rect 159326 16718 159562 16954
rect 159646 16718 159882 16954
rect 159326 16398 159562 16634
rect 159646 16398 159882 16634
rect 159326 -3462 159562 -3226
rect 159646 -3462 159882 -3226
rect 159326 -3782 159562 -3546
rect 159646 -3782 159882 -3546
rect 163826 489218 164062 489454
rect 164146 489218 164382 489454
rect 163826 488898 164062 489134
rect 164146 488898 164382 489134
rect 163826 453218 164062 453454
rect 164146 453218 164382 453454
rect 163826 452898 164062 453134
rect 164146 452898 164382 453134
rect 163826 417218 164062 417454
rect 164146 417218 164382 417454
rect 163826 416898 164062 417134
rect 164146 416898 164382 417134
rect 163826 381218 164062 381454
rect 164146 381218 164382 381454
rect 163826 380898 164062 381134
rect 164146 380898 164382 381134
rect 163826 345218 164062 345454
rect 164146 345218 164382 345454
rect 163826 344898 164062 345134
rect 164146 344898 164382 345134
rect 163826 309218 164062 309454
rect 164146 309218 164382 309454
rect 163826 308898 164062 309134
rect 164146 308898 164382 309134
rect 163826 273218 164062 273454
rect 164146 273218 164382 273454
rect 163826 272898 164062 273134
rect 164146 272898 164382 273134
rect 163826 237218 164062 237454
rect 164146 237218 164382 237454
rect 163826 236898 164062 237134
rect 164146 236898 164382 237134
rect 163826 201218 164062 201454
rect 164146 201218 164382 201454
rect 163826 200898 164062 201134
rect 164146 200898 164382 201134
rect 163826 165218 164062 165454
rect 164146 165218 164382 165454
rect 163826 164898 164062 165134
rect 164146 164898 164382 165134
rect 163826 129218 164062 129454
rect 164146 129218 164382 129454
rect 163826 128898 164062 129134
rect 164146 128898 164382 129134
rect 163826 93218 164062 93454
rect 164146 93218 164382 93454
rect 163826 92898 164062 93134
rect 164146 92898 164382 93134
rect 163826 57218 164062 57454
rect 164146 57218 164382 57454
rect 163826 56898 164062 57134
rect 164146 56898 164382 57134
rect 163826 21218 164062 21454
rect 164146 21218 164382 21454
rect 163826 20898 164062 21134
rect 164146 20898 164382 21134
rect 163826 -4422 164062 -4186
rect 164146 -4422 164382 -4186
rect 163826 -4742 164062 -4506
rect 164146 -4742 164382 -4506
rect 168326 493718 168562 493954
rect 168646 493718 168882 493954
rect 168326 493398 168562 493634
rect 168646 493398 168882 493634
rect 168326 457718 168562 457954
rect 168646 457718 168882 457954
rect 168326 457398 168562 457634
rect 168646 457398 168882 457634
rect 168326 421718 168562 421954
rect 168646 421718 168882 421954
rect 168326 421398 168562 421634
rect 168646 421398 168882 421634
rect 168326 385718 168562 385954
rect 168646 385718 168882 385954
rect 168326 385398 168562 385634
rect 168646 385398 168882 385634
rect 168326 349718 168562 349954
rect 168646 349718 168882 349954
rect 168326 349398 168562 349634
rect 168646 349398 168882 349634
rect 168326 313718 168562 313954
rect 168646 313718 168882 313954
rect 168326 313398 168562 313634
rect 168646 313398 168882 313634
rect 168326 277718 168562 277954
rect 168646 277718 168882 277954
rect 168326 277398 168562 277634
rect 168646 277398 168882 277634
rect 168326 241718 168562 241954
rect 168646 241718 168882 241954
rect 168326 241398 168562 241634
rect 168646 241398 168882 241634
rect 168326 205718 168562 205954
rect 168646 205718 168882 205954
rect 168326 205398 168562 205634
rect 168646 205398 168882 205634
rect 168326 169718 168562 169954
rect 168646 169718 168882 169954
rect 168326 169398 168562 169634
rect 168646 169398 168882 169634
rect 168326 133718 168562 133954
rect 168646 133718 168882 133954
rect 168326 133398 168562 133634
rect 168646 133398 168882 133634
rect 168326 97718 168562 97954
rect 168646 97718 168882 97954
rect 168326 97398 168562 97634
rect 168646 97398 168882 97634
rect 168326 61718 168562 61954
rect 168646 61718 168882 61954
rect 168326 61398 168562 61634
rect 168646 61398 168882 61634
rect 168326 25718 168562 25954
rect 168646 25718 168882 25954
rect 168326 25398 168562 25634
rect 168646 25398 168882 25634
rect 168326 -5382 168562 -5146
rect 168646 -5382 168882 -5146
rect 168326 -5702 168562 -5466
rect 168646 -5702 168882 -5466
rect 172826 462218 173062 462454
rect 173146 462218 173382 462454
rect 172826 461898 173062 462134
rect 173146 461898 173382 462134
rect 172826 426218 173062 426454
rect 173146 426218 173382 426454
rect 172826 425898 173062 426134
rect 173146 425898 173382 426134
rect 172826 390218 173062 390454
rect 173146 390218 173382 390454
rect 172826 389898 173062 390134
rect 173146 389898 173382 390134
rect 172826 354218 173062 354454
rect 173146 354218 173382 354454
rect 172826 353898 173062 354134
rect 173146 353898 173382 354134
rect 172826 318218 173062 318454
rect 173146 318218 173382 318454
rect 172826 317898 173062 318134
rect 173146 317898 173382 318134
rect 172826 282218 173062 282454
rect 173146 282218 173382 282454
rect 172826 281898 173062 282134
rect 173146 281898 173382 282134
rect 172826 246218 173062 246454
rect 173146 246218 173382 246454
rect 172826 245898 173062 246134
rect 173146 245898 173382 246134
rect 172826 210218 173062 210454
rect 173146 210218 173382 210454
rect 172826 209898 173062 210134
rect 173146 209898 173382 210134
rect 172826 174218 173062 174454
rect 173146 174218 173382 174454
rect 172826 173898 173062 174134
rect 173146 173898 173382 174134
rect 172826 138218 173062 138454
rect 173146 138218 173382 138454
rect 172826 137898 173062 138134
rect 173146 137898 173382 138134
rect 172826 102218 173062 102454
rect 173146 102218 173382 102454
rect 172826 101898 173062 102134
rect 173146 101898 173382 102134
rect 172826 66218 173062 66454
rect 173146 66218 173382 66454
rect 172826 65898 173062 66134
rect 173146 65898 173382 66134
rect 172826 30218 173062 30454
rect 173146 30218 173382 30454
rect 172826 29898 173062 30134
rect 173146 29898 173382 30134
rect 172826 -6342 173062 -6106
rect 173146 -6342 173382 -6106
rect 172826 -6662 173062 -6426
rect 173146 -6662 173382 -6426
rect 177326 466718 177562 466954
rect 177646 466718 177882 466954
rect 177326 466398 177562 466634
rect 177646 466398 177882 466634
rect 177326 430718 177562 430954
rect 177646 430718 177882 430954
rect 177326 430398 177562 430634
rect 177646 430398 177882 430634
rect 177326 394718 177562 394954
rect 177646 394718 177882 394954
rect 177326 394398 177562 394634
rect 177646 394398 177882 394634
rect 177326 358718 177562 358954
rect 177646 358718 177882 358954
rect 177326 358398 177562 358634
rect 177646 358398 177882 358634
rect 177326 322718 177562 322954
rect 177646 322718 177882 322954
rect 177326 322398 177562 322634
rect 177646 322398 177882 322634
rect 177326 286718 177562 286954
rect 177646 286718 177882 286954
rect 177326 286398 177562 286634
rect 177646 286398 177882 286634
rect 177326 250718 177562 250954
rect 177646 250718 177882 250954
rect 177326 250398 177562 250634
rect 177646 250398 177882 250634
rect 177326 214718 177562 214954
rect 177646 214718 177882 214954
rect 177326 214398 177562 214634
rect 177646 214398 177882 214634
rect 177326 178718 177562 178954
rect 177646 178718 177882 178954
rect 177326 178398 177562 178634
rect 177646 178398 177882 178634
rect 177326 142718 177562 142954
rect 177646 142718 177882 142954
rect 177326 142398 177562 142634
rect 177646 142398 177882 142634
rect 177326 106718 177562 106954
rect 177646 106718 177882 106954
rect 177326 106398 177562 106634
rect 177646 106398 177882 106634
rect 177326 70718 177562 70954
rect 177646 70718 177882 70954
rect 177326 70398 177562 70634
rect 177646 70398 177882 70634
rect 177326 34718 177562 34954
rect 177646 34718 177882 34954
rect 177326 34398 177562 34634
rect 177646 34398 177882 34634
rect 177326 -7302 177562 -7066
rect 177646 -7302 177882 -7066
rect 177326 -7622 177562 -7386
rect 177646 -7622 177882 -7386
rect 181826 471218 182062 471454
rect 182146 471218 182382 471454
rect 181826 470898 182062 471134
rect 182146 470898 182382 471134
rect 181826 435218 182062 435454
rect 182146 435218 182382 435454
rect 181826 434898 182062 435134
rect 182146 434898 182382 435134
rect 181826 399218 182062 399454
rect 182146 399218 182382 399454
rect 181826 398898 182062 399134
rect 182146 398898 182382 399134
rect 181826 363218 182062 363454
rect 182146 363218 182382 363454
rect 181826 362898 182062 363134
rect 182146 362898 182382 363134
rect 181826 327218 182062 327454
rect 182146 327218 182382 327454
rect 181826 326898 182062 327134
rect 182146 326898 182382 327134
rect 181826 291218 182062 291454
rect 182146 291218 182382 291454
rect 181826 290898 182062 291134
rect 182146 290898 182382 291134
rect 181826 255218 182062 255454
rect 182146 255218 182382 255454
rect 181826 254898 182062 255134
rect 182146 254898 182382 255134
rect 181826 219218 182062 219454
rect 182146 219218 182382 219454
rect 181826 218898 182062 219134
rect 182146 218898 182382 219134
rect 181826 183218 182062 183454
rect 182146 183218 182382 183454
rect 181826 182898 182062 183134
rect 182146 182898 182382 183134
rect 181826 147218 182062 147454
rect 182146 147218 182382 147454
rect 181826 146898 182062 147134
rect 182146 146898 182382 147134
rect 181826 111218 182062 111454
rect 182146 111218 182382 111454
rect 181826 110898 182062 111134
rect 182146 110898 182382 111134
rect 181826 75218 182062 75454
rect 182146 75218 182382 75454
rect 181826 74898 182062 75134
rect 182146 74898 182382 75134
rect 181826 39218 182062 39454
rect 182146 39218 182382 39454
rect 181826 38898 182062 39134
rect 182146 38898 182382 39134
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 186326 475718 186562 475954
rect 186646 475718 186882 475954
rect 186326 475398 186562 475634
rect 186646 475398 186882 475634
rect 186326 439718 186562 439954
rect 186646 439718 186882 439954
rect 186326 439398 186562 439634
rect 186646 439398 186882 439634
rect 186326 403718 186562 403954
rect 186646 403718 186882 403954
rect 186326 403398 186562 403634
rect 186646 403398 186882 403634
rect 186326 367718 186562 367954
rect 186646 367718 186882 367954
rect 186326 367398 186562 367634
rect 186646 367398 186882 367634
rect 186326 331718 186562 331954
rect 186646 331718 186882 331954
rect 186326 331398 186562 331634
rect 186646 331398 186882 331634
rect 186326 295718 186562 295954
rect 186646 295718 186882 295954
rect 186326 295398 186562 295634
rect 186646 295398 186882 295634
rect 186326 259718 186562 259954
rect 186646 259718 186882 259954
rect 186326 259398 186562 259634
rect 186646 259398 186882 259634
rect 186326 223718 186562 223954
rect 186646 223718 186882 223954
rect 186326 223398 186562 223634
rect 186646 223398 186882 223634
rect 186326 187718 186562 187954
rect 186646 187718 186882 187954
rect 186326 187398 186562 187634
rect 186646 187398 186882 187634
rect 186326 151718 186562 151954
rect 186646 151718 186882 151954
rect 186326 151398 186562 151634
rect 186646 151398 186882 151634
rect 186326 115718 186562 115954
rect 186646 115718 186882 115954
rect 186326 115398 186562 115634
rect 186646 115398 186882 115634
rect 186326 79718 186562 79954
rect 186646 79718 186882 79954
rect 186326 79398 186562 79634
rect 186646 79398 186882 79634
rect 186326 43718 186562 43954
rect 186646 43718 186882 43954
rect 186326 43398 186562 43634
rect 186646 43398 186882 43634
rect 186326 7718 186562 7954
rect 186646 7718 186882 7954
rect 186326 7398 186562 7634
rect 186646 7398 186882 7634
rect 186326 -1542 186562 -1306
rect 186646 -1542 186882 -1306
rect 186326 -1862 186562 -1626
rect 186646 -1862 186882 -1626
rect 190826 480218 191062 480454
rect 191146 480218 191382 480454
rect 190826 479898 191062 480134
rect 191146 479898 191382 480134
rect 190826 444218 191062 444454
rect 191146 444218 191382 444454
rect 190826 443898 191062 444134
rect 191146 443898 191382 444134
rect 190826 408218 191062 408454
rect 191146 408218 191382 408454
rect 190826 407898 191062 408134
rect 191146 407898 191382 408134
rect 190826 372218 191062 372454
rect 191146 372218 191382 372454
rect 190826 371898 191062 372134
rect 191146 371898 191382 372134
rect 190826 336218 191062 336454
rect 191146 336218 191382 336454
rect 190826 335898 191062 336134
rect 191146 335898 191382 336134
rect 190826 300218 191062 300454
rect 191146 300218 191382 300454
rect 190826 299898 191062 300134
rect 191146 299898 191382 300134
rect 190826 264218 191062 264454
rect 191146 264218 191382 264454
rect 190826 263898 191062 264134
rect 191146 263898 191382 264134
rect 190826 228218 191062 228454
rect 191146 228218 191382 228454
rect 190826 227898 191062 228134
rect 191146 227898 191382 228134
rect 190826 192218 191062 192454
rect 191146 192218 191382 192454
rect 190826 191898 191062 192134
rect 191146 191898 191382 192134
rect 190826 156218 191062 156454
rect 191146 156218 191382 156454
rect 190826 155898 191062 156134
rect 191146 155898 191382 156134
rect 190826 120218 191062 120454
rect 191146 120218 191382 120454
rect 190826 119898 191062 120134
rect 191146 119898 191382 120134
rect 190826 84218 191062 84454
rect 191146 84218 191382 84454
rect 190826 83898 191062 84134
rect 191146 83898 191382 84134
rect 190826 48218 191062 48454
rect 191146 48218 191382 48454
rect 190826 47898 191062 48134
rect 191146 47898 191382 48134
rect 190826 12218 191062 12454
rect 191146 12218 191382 12454
rect 190826 11898 191062 12134
rect 191146 11898 191382 12134
rect 190826 -2502 191062 -2266
rect 191146 -2502 191382 -2266
rect 190826 -2822 191062 -2586
rect 191146 -2822 191382 -2586
rect 195326 484718 195562 484954
rect 195646 484718 195882 484954
rect 195326 484398 195562 484634
rect 195646 484398 195882 484634
rect 195326 448718 195562 448954
rect 195646 448718 195882 448954
rect 195326 448398 195562 448634
rect 195646 448398 195882 448634
rect 195326 412718 195562 412954
rect 195646 412718 195882 412954
rect 195326 412398 195562 412634
rect 195646 412398 195882 412634
rect 195326 376718 195562 376954
rect 195646 376718 195882 376954
rect 195326 376398 195562 376634
rect 195646 376398 195882 376634
rect 195326 340718 195562 340954
rect 195646 340718 195882 340954
rect 195326 340398 195562 340634
rect 195646 340398 195882 340634
rect 195326 304718 195562 304954
rect 195646 304718 195882 304954
rect 195326 304398 195562 304634
rect 195646 304398 195882 304634
rect 195326 268718 195562 268954
rect 195646 268718 195882 268954
rect 195326 268398 195562 268634
rect 195646 268398 195882 268634
rect 195326 232718 195562 232954
rect 195646 232718 195882 232954
rect 195326 232398 195562 232634
rect 195646 232398 195882 232634
rect 195326 196718 195562 196954
rect 195646 196718 195882 196954
rect 195326 196398 195562 196634
rect 195646 196398 195882 196634
rect 195326 160718 195562 160954
rect 195646 160718 195882 160954
rect 195326 160398 195562 160634
rect 195646 160398 195882 160634
rect 195326 124718 195562 124954
rect 195646 124718 195882 124954
rect 195326 124398 195562 124634
rect 195646 124398 195882 124634
rect 195326 88718 195562 88954
rect 195646 88718 195882 88954
rect 195326 88398 195562 88634
rect 195646 88398 195882 88634
rect 195326 52718 195562 52954
rect 195646 52718 195882 52954
rect 195326 52398 195562 52634
rect 195646 52398 195882 52634
rect 195326 16718 195562 16954
rect 195646 16718 195882 16954
rect 195326 16398 195562 16634
rect 195646 16398 195882 16634
rect 195326 -3462 195562 -3226
rect 195646 -3462 195882 -3226
rect 195326 -3782 195562 -3546
rect 195646 -3782 195882 -3546
rect 199826 708442 200062 708678
rect 200146 708442 200382 708678
rect 199826 708122 200062 708358
rect 200146 708122 200382 708358
rect 199826 669218 200062 669454
rect 200146 669218 200382 669454
rect 199826 668898 200062 669134
rect 200146 668898 200382 669134
rect 199826 633218 200062 633454
rect 200146 633218 200382 633454
rect 199826 632898 200062 633134
rect 200146 632898 200382 633134
rect 199826 597218 200062 597454
rect 200146 597218 200382 597454
rect 199826 596898 200062 597134
rect 200146 596898 200382 597134
rect 199826 561218 200062 561454
rect 200146 561218 200382 561454
rect 199826 560898 200062 561134
rect 200146 560898 200382 561134
rect 199826 525218 200062 525454
rect 200146 525218 200382 525454
rect 199826 524898 200062 525134
rect 200146 524898 200382 525134
rect 199826 489218 200062 489454
rect 200146 489218 200382 489454
rect 199826 488898 200062 489134
rect 200146 488898 200382 489134
rect 199826 453218 200062 453454
rect 200146 453218 200382 453454
rect 199826 452898 200062 453134
rect 200146 452898 200382 453134
rect 199826 417218 200062 417454
rect 200146 417218 200382 417454
rect 199826 416898 200062 417134
rect 200146 416898 200382 417134
rect 199826 381218 200062 381454
rect 200146 381218 200382 381454
rect 199826 380898 200062 381134
rect 200146 380898 200382 381134
rect 199826 345218 200062 345454
rect 200146 345218 200382 345454
rect 199826 344898 200062 345134
rect 200146 344898 200382 345134
rect 199826 309218 200062 309454
rect 200146 309218 200382 309454
rect 199826 308898 200062 309134
rect 200146 308898 200382 309134
rect 199826 273218 200062 273454
rect 200146 273218 200382 273454
rect 199826 272898 200062 273134
rect 200146 272898 200382 273134
rect 199826 237218 200062 237454
rect 200146 237218 200382 237454
rect 199826 236898 200062 237134
rect 200146 236898 200382 237134
rect 199826 201218 200062 201454
rect 200146 201218 200382 201454
rect 199826 200898 200062 201134
rect 200146 200898 200382 201134
rect 199826 165218 200062 165454
rect 200146 165218 200382 165454
rect 199826 164898 200062 165134
rect 200146 164898 200382 165134
rect 199826 129218 200062 129454
rect 200146 129218 200382 129454
rect 199826 128898 200062 129134
rect 200146 128898 200382 129134
rect 199826 93218 200062 93454
rect 200146 93218 200382 93454
rect 199826 92898 200062 93134
rect 200146 92898 200382 93134
rect 199826 57218 200062 57454
rect 200146 57218 200382 57454
rect 199826 56898 200062 57134
rect 200146 56898 200382 57134
rect 199826 21218 200062 21454
rect 200146 21218 200382 21454
rect 199826 20898 200062 21134
rect 200146 20898 200382 21134
rect 199826 -4422 200062 -4186
rect 200146 -4422 200382 -4186
rect 199826 -4742 200062 -4506
rect 200146 -4742 200382 -4506
rect 204326 709402 204562 709638
rect 204646 709402 204882 709638
rect 204326 709082 204562 709318
rect 204646 709082 204882 709318
rect 204326 673718 204562 673954
rect 204646 673718 204882 673954
rect 204326 673398 204562 673634
rect 204646 673398 204882 673634
rect 204326 637718 204562 637954
rect 204646 637718 204882 637954
rect 204326 637398 204562 637634
rect 204646 637398 204882 637634
rect 204326 601718 204562 601954
rect 204646 601718 204882 601954
rect 204326 601398 204562 601634
rect 204646 601398 204882 601634
rect 204326 565718 204562 565954
rect 204646 565718 204882 565954
rect 204326 565398 204562 565634
rect 204646 565398 204882 565634
rect 204326 529718 204562 529954
rect 204646 529718 204882 529954
rect 204326 529398 204562 529634
rect 204646 529398 204882 529634
rect 204326 493718 204562 493954
rect 204646 493718 204882 493954
rect 204326 493398 204562 493634
rect 204646 493398 204882 493634
rect 204326 457718 204562 457954
rect 204646 457718 204882 457954
rect 204326 457398 204562 457634
rect 204646 457398 204882 457634
rect 204326 421718 204562 421954
rect 204646 421718 204882 421954
rect 204326 421398 204562 421634
rect 204646 421398 204882 421634
rect 204326 385718 204562 385954
rect 204646 385718 204882 385954
rect 204326 385398 204562 385634
rect 204646 385398 204882 385634
rect 204326 349718 204562 349954
rect 204646 349718 204882 349954
rect 204326 349398 204562 349634
rect 204646 349398 204882 349634
rect 204326 313718 204562 313954
rect 204646 313718 204882 313954
rect 204326 313398 204562 313634
rect 204646 313398 204882 313634
rect 204326 277718 204562 277954
rect 204646 277718 204882 277954
rect 204326 277398 204562 277634
rect 204646 277398 204882 277634
rect 204326 241718 204562 241954
rect 204646 241718 204882 241954
rect 204326 241398 204562 241634
rect 204646 241398 204882 241634
rect 204326 205718 204562 205954
rect 204646 205718 204882 205954
rect 204326 205398 204562 205634
rect 204646 205398 204882 205634
rect 204326 169718 204562 169954
rect 204646 169718 204882 169954
rect 204326 169398 204562 169634
rect 204646 169398 204882 169634
rect 204326 133718 204562 133954
rect 204646 133718 204882 133954
rect 204326 133398 204562 133634
rect 204646 133398 204882 133634
rect 204326 97718 204562 97954
rect 204646 97718 204882 97954
rect 204326 97398 204562 97634
rect 204646 97398 204882 97634
rect 204326 61718 204562 61954
rect 204646 61718 204882 61954
rect 204326 61398 204562 61634
rect 204646 61398 204882 61634
rect 204326 25718 204562 25954
rect 204646 25718 204882 25954
rect 204326 25398 204562 25634
rect 204646 25398 204882 25634
rect 204326 -5382 204562 -5146
rect 204646 -5382 204882 -5146
rect 204326 -5702 204562 -5466
rect 204646 -5702 204882 -5466
rect 208826 710362 209062 710598
rect 209146 710362 209382 710598
rect 208826 710042 209062 710278
rect 209146 710042 209382 710278
rect 208826 678218 209062 678454
rect 209146 678218 209382 678454
rect 208826 677898 209062 678134
rect 209146 677898 209382 678134
rect 208826 642218 209062 642454
rect 209146 642218 209382 642454
rect 208826 641898 209062 642134
rect 209146 641898 209382 642134
rect 208826 606218 209062 606454
rect 209146 606218 209382 606454
rect 208826 605898 209062 606134
rect 209146 605898 209382 606134
rect 208826 570218 209062 570454
rect 209146 570218 209382 570454
rect 208826 569898 209062 570134
rect 209146 569898 209382 570134
rect 208826 534218 209062 534454
rect 209146 534218 209382 534454
rect 208826 533898 209062 534134
rect 209146 533898 209382 534134
rect 208826 498218 209062 498454
rect 209146 498218 209382 498454
rect 208826 497898 209062 498134
rect 209146 497898 209382 498134
rect 208826 462218 209062 462454
rect 209146 462218 209382 462454
rect 208826 461898 209062 462134
rect 209146 461898 209382 462134
rect 208826 426218 209062 426454
rect 209146 426218 209382 426454
rect 208826 425898 209062 426134
rect 209146 425898 209382 426134
rect 208826 390218 209062 390454
rect 209146 390218 209382 390454
rect 208826 389898 209062 390134
rect 209146 389898 209382 390134
rect 208826 354218 209062 354454
rect 209146 354218 209382 354454
rect 208826 353898 209062 354134
rect 209146 353898 209382 354134
rect 208826 318218 209062 318454
rect 209146 318218 209382 318454
rect 208826 317898 209062 318134
rect 209146 317898 209382 318134
rect 208826 282218 209062 282454
rect 209146 282218 209382 282454
rect 208826 281898 209062 282134
rect 209146 281898 209382 282134
rect 208826 246218 209062 246454
rect 209146 246218 209382 246454
rect 208826 245898 209062 246134
rect 209146 245898 209382 246134
rect 208826 210218 209062 210454
rect 209146 210218 209382 210454
rect 208826 209898 209062 210134
rect 209146 209898 209382 210134
rect 208826 174218 209062 174454
rect 209146 174218 209382 174454
rect 208826 173898 209062 174134
rect 209146 173898 209382 174134
rect 208826 138218 209062 138454
rect 209146 138218 209382 138454
rect 208826 137898 209062 138134
rect 209146 137898 209382 138134
rect 208826 102218 209062 102454
rect 209146 102218 209382 102454
rect 208826 101898 209062 102134
rect 209146 101898 209382 102134
rect 208826 66218 209062 66454
rect 209146 66218 209382 66454
rect 208826 65898 209062 66134
rect 209146 65898 209382 66134
rect 208826 30218 209062 30454
rect 209146 30218 209382 30454
rect 208826 29898 209062 30134
rect 209146 29898 209382 30134
rect 208826 -6342 209062 -6106
rect 209146 -6342 209382 -6106
rect 208826 -6662 209062 -6426
rect 209146 -6662 209382 -6426
rect 213326 711322 213562 711558
rect 213646 711322 213882 711558
rect 213326 711002 213562 711238
rect 213646 711002 213882 711238
rect 213326 682718 213562 682954
rect 213646 682718 213882 682954
rect 213326 682398 213562 682634
rect 213646 682398 213882 682634
rect 213326 646718 213562 646954
rect 213646 646718 213882 646954
rect 213326 646398 213562 646634
rect 213646 646398 213882 646634
rect 213326 610718 213562 610954
rect 213646 610718 213882 610954
rect 213326 610398 213562 610634
rect 213646 610398 213882 610634
rect 213326 574718 213562 574954
rect 213646 574718 213882 574954
rect 213326 574398 213562 574634
rect 213646 574398 213882 574634
rect 213326 538718 213562 538954
rect 213646 538718 213882 538954
rect 213326 538398 213562 538634
rect 213646 538398 213882 538634
rect 213326 502718 213562 502954
rect 213646 502718 213882 502954
rect 213326 502398 213562 502634
rect 213646 502398 213882 502634
rect 213326 466718 213562 466954
rect 213646 466718 213882 466954
rect 213326 466398 213562 466634
rect 213646 466398 213882 466634
rect 213326 430718 213562 430954
rect 213646 430718 213882 430954
rect 213326 430398 213562 430634
rect 213646 430398 213882 430634
rect 213326 394718 213562 394954
rect 213646 394718 213882 394954
rect 213326 394398 213562 394634
rect 213646 394398 213882 394634
rect 213326 358718 213562 358954
rect 213646 358718 213882 358954
rect 213326 358398 213562 358634
rect 213646 358398 213882 358634
rect 213326 322718 213562 322954
rect 213646 322718 213882 322954
rect 213326 322398 213562 322634
rect 213646 322398 213882 322634
rect 213326 286718 213562 286954
rect 213646 286718 213882 286954
rect 213326 286398 213562 286634
rect 213646 286398 213882 286634
rect 213326 250718 213562 250954
rect 213646 250718 213882 250954
rect 213326 250398 213562 250634
rect 213646 250398 213882 250634
rect 213326 214718 213562 214954
rect 213646 214718 213882 214954
rect 213326 214398 213562 214634
rect 213646 214398 213882 214634
rect 213326 178718 213562 178954
rect 213646 178718 213882 178954
rect 213326 178398 213562 178634
rect 213646 178398 213882 178634
rect 213326 142718 213562 142954
rect 213646 142718 213882 142954
rect 213326 142398 213562 142634
rect 213646 142398 213882 142634
rect 213326 106718 213562 106954
rect 213646 106718 213882 106954
rect 213326 106398 213562 106634
rect 213646 106398 213882 106634
rect 213326 70718 213562 70954
rect 213646 70718 213882 70954
rect 213326 70398 213562 70634
rect 213646 70398 213882 70634
rect 213326 34718 213562 34954
rect 213646 34718 213882 34954
rect 213326 34398 213562 34634
rect 213646 34398 213882 34634
rect 213326 -7302 213562 -7066
rect 213646 -7302 213882 -7066
rect 213326 -7622 213562 -7386
rect 213646 -7622 213882 -7386
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 217826 651218 218062 651454
rect 218146 651218 218382 651454
rect 217826 650898 218062 651134
rect 218146 650898 218382 651134
rect 217826 615218 218062 615454
rect 218146 615218 218382 615454
rect 217826 614898 218062 615134
rect 218146 614898 218382 615134
rect 217826 579218 218062 579454
rect 218146 579218 218382 579454
rect 217826 578898 218062 579134
rect 218146 578898 218382 579134
rect 217826 543218 218062 543454
rect 218146 543218 218382 543454
rect 217826 542898 218062 543134
rect 218146 542898 218382 543134
rect 217826 507218 218062 507454
rect 218146 507218 218382 507454
rect 217826 506898 218062 507134
rect 218146 506898 218382 507134
rect 217826 471218 218062 471454
rect 218146 471218 218382 471454
rect 217826 470898 218062 471134
rect 218146 470898 218382 471134
rect 217826 435218 218062 435454
rect 218146 435218 218382 435454
rect 217826 434898 218062 435134
rect 218146 434898 218382 435134
rect 217826 399218 218062 399454
rect 218146 399218 218382 399454
rect 217826 398898 218062 399134
rect 218146 398898 218382 399134
rect 217826 363218 218062 363454
rect 218146 363218 218382 363454
rect 217826 362898 218062 363134
rect 218146 362898 218382 363134
rect 217826 327218 218062 327454
rect 218146 327218 218382 327454
rect 217826 326898 218062 327134
rect 218146 326898 218382 327134
rect 217826 291218 218062 291454
rect 218146 291218 218382 291454
rect 217826 290898 218062 291134
rect 218146 290898 218382 291134
rect 217826 255218 218062 255454
rect 218146 255218 218382 255454
rect 217826 254898 218062 255134
rect 218146 254898 218382 255134
rect 217826 219218 218062 219454
rect 218146 219218 218382 219454
rect 217826 218898 218062 219134
rect 218146 218898 218382 219134
rect 217826 183218 218062 183454
rect 218146 183218 218382 183454
rect 217826 182898 218062 183134
rect 218146 182898 218382 183134
rect 217826 147218 218062 147454
rect 218146 147218 218382 147454
rect 217826 146898 218062 147134
rect 218146 146898 218382 147134
rect 217826 111218 218062 111454
rect 218146 111218 218382 111454
rect 217826 110898 218062 111134
rect 218146 110898 218382 111134
rect 217826 75218 218062 75454
rect 218146 75218 218382 75454
rect 217826 74898 218062 75134
rect 218146 74898 218382 75134
rect 217826 39218 218062 39454
rect 218146 39218 218382 39454
rect 217826 38898 218062 39134
rect 218146 38898 218382 39134
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 222326 705562 222562 705798
rect 222646 705562 222882 705798
rect 222326 705242 222562 705478
rect 222646 705242 222882 705478
rect 222326 691718 222562 691954
rect 222646 691718 222882 691954
rect 222326 691398 222562 691634
rect 222646 691398 222882 691634
rect 222326 655718 222562 655954
rect 222646 655718 222882 655954
rect 222326 655398 222562 655634
rect 222646 655398 222882 655634
rect 222326 619718 222562 619954
rect 222646 619718 222882 619954
rect 222326 619398 222562 619634
rect 222646 619398 222882 619634
rect 222326 583718 222562 583954
rect 222646 583718 222882 583954
rect 222326 583398 222562 583634
rect 222646 583398 222882 583634
rect 222326 547718 222562 547954
rect 222646 547718 222882 547954
rect 222326 547398 222562 547634
rect 222646 547398 222882 547634
rect 222326 511718 222562 511954
rect 222646 511718 222882 511954
rect 222326 511398 222562 511634
rect 222646 511398 222882 511634
rect 222326 475718 222562 475954
rect 222646 475718 222882 475954
rect 222326 475398 222562 475634
rect 222646 475398 222882 475634
rect 222326 439718 222562 439954
rect 222646 439718 222882 439954
rect 222326 439398 222562 439634
rect 222646 439398 222882 439634
rect 222326 403718 222562 403954
rect 222646 403718 222882 403954
rect 222326 403398 222562 403634
rect 222646 403398 222882 403634
rect 222326 367718 222562 367954
rect 222646 367718 222882 367954
rect 222326 367398 222562 367634
rect 222646 367398 222882 367634
rect 222326 331718 222562 331954
rect 222646 331718 222882 331954
rect 222326 331398 222562 331634
rect 222646 331398 222882 331634
rect 222326 295718 222562 295954
rect 222646 295718 222882 295954
rect 222326 295398 222562 295634
rect 222646 295398 222882 295634
rect 222326 259718 222562 259954
rect 222646 259718 222882 259954
rect 222326 259398 222562 259634
rect 222646 259398 222882 259634
rect 222326 223718 222562 223954
rect 222646 223718 222882 223954
rect 222326 223398 222562 223634
rect 222646 223398 222882 223634
rect 222326 187718 222562 187954
rect 222646 187718 222882 187954
rect 222326 187398 222562 187634
rect 222646 187398 222882 187634
rect 222326 151718 222562 151954
rect 222646 151718 222882 151954
rect 222326 151398 222562 151634
rect 222646 151398 222882 151634
rect 222326 115718 222562 115954
rect 222646 115718 222882 115954
rect 222326 115398 222562 115634
rect 222646 115398 222882 115634
rect 222326 79718 222562 79954
rect 222646 79718 222882 79954
rect 222326 79398 222562 79634
rect 222646 79398 222882 79634
rect 222326 43718 222562 43954
rect 222646 43718 222882 43954
rect 222326 43398 222562 43634
rect 222646 43398 222882 43634
rect 222326 7718 222562 7954
rect 222646 7718 222882 7954
rect 222326 7398 222562 7634
rect 222646 7398 222882 7634
rect 222326 -1542 222562 -1306
rect 222646 -1542 222882 -1306
rect 222326 -1862 222562 -1626
rect 222646 -1862 222882 -1626
rect 226826 706522 227062 706758
rect 227146 706522 227382 706758
rect 226826 706202 227062 706438
rect 227146 706202 227382 706438
rect 226826 696218 227062 696454
rect 227146 696218 227382 696454
rect 226826 695898 227062 696134
rect 227146 695898 227382 696134
rect 226826 660218 227062 660454
rect 227146 660218 227382 660454
rect 226826 659898 227062 660134
rect 227146 659898 227382 660134
rect 226826 624218 227062 624454
rect 227146 624218 227382 624454
rect 226826 623898 227062 624134
rect 227146 623898 227382 624134
rect 226826 588218 227062 588454
rect 227146 588218 227382 588454
rect 226826 587898 227062 588134
rect 227146 587898 227382 588134
rect 226826 552218 227062 552454
rect 227146 552218 227382 552454
rect 226826 551898 227062 552134
rect 227146 551898 227382 552134
rect 226826 516218 227062 516454
rect 227146 516218 227382 516454
rect 226826 515898 227062 516134
rect 227146 515898 227382 516134
rect 226826 480218 227062 480454
rect 227146 480218 227382 480454
rect 226826 479898 227062 480134
rect 227146 479898 227382 480134
rect 226826 444218 227062 444454
rect 227146 444218 227382 444454
rect 226826 443898 227062 444134
rect 227146 443898 227382 444134
rect 226826 408218 227062 408454
rect 227146 408218 227382 408454
rect 226826 407898 227062 408134
rect 227146 407898 227382 408134
rect 226826 372218 227062 372454
rect 227146 372218 227382 372454
rect 226826 371898 227062 372134
rect 227146 371898 227382 372134
rect 226826 336218 227062 336454
rect 227146 336218 227382 336454
rect 226826 335898 227062 336134
rect 227146 335898 227382 336134
rect 226826 300218 227062 300454
rect 227146 300218 227382 300454
rect 226826 299898 227062 300134
rect 227146 299898 227382 300134
rect 226826 264218 227062 264454
rect 227146 264218 227382 264454
rect 226826 263898 227062 264134
rect 227146 263898 227382 264134
rect 226826 228218 227062 228454
rect 227146 228218 227382 228454
rect 226826 227898 227062 228134
rect 227146 227898 227382 228134
rect 226826 192218 227062 192454
rect 227146 192218 227382 192454
rect 226826 191898 227062 192134
rect 227146 191898 227382 192134
rect 226826 156218 227062 156454
rect 227146 156218 227382 156454
rect 226826 155898 227062 156134
rect 227146 155898 227382 156134
rect 226826 120218 227062 120454
rect 227146 120218 227382 120454
rect 226826 119898 227062 120134
rect 227146 119898 227382 120134
rect 226826 84218 227062 84454
rect 227146 84218 227382 84454
rect 226826 83898 227062 84134
rect 227146 83898 227382 84134
rect 226826 48218 227062 48454
rect 227146 48218 227382 48454
rect 226826 47898 227062 48134
rect 227146 47898 227382 48134
rect 226826 12218 227062 12454
rect 227146 12218 227382 12454
rect 226826 11898 227062 12134
rect 227146 11898 227382 12134
rect 226826 -2502 227062 -2266
rect 227146 -2502 227382 -2266
rect 226826 -2822 227062 -2586
rect 227146 -2822 227382 -2586
rect 231326 707482 231562 707718
rect 231646 707482 231882 707718
rect 231326 707162 231562 707398
rect 231646 707162 231882 707398
rect 231326 700718 231562 700954
rect 231646 700718 231882 700954
rect 231326 700398 231562 700634
rect 231646 700398 231882 700634
rect 231326 664718 231562 664954
rect 231646 664718 231882 664954
rect 231326 664398 231562 664634
rect 231646 664398 231882 664634
rect 231326 628718 231562 628954
rect 231646 628718 231882 628954
rect 231326 628398 231562 628634
rect 231646 628398 231882 628634
rect 231326 592718 231562 592954
rect 231646 592718 231882 592954
rect 231326 592398 231562 592634
rect 231646 592398 231882 592634
rect 231326 556718 231562 556954
rect 231646 556718 231882 556954
rect 231326 556398 231562 556634
rect 231646 556398 231882 556634
rect 231326 520718 231562 520954
rect 231646 520718 231882 520954
rect 231326 520398 231562 520634
rect 231646 520398 231882 520634
rect 231326 484718 231562 484954
rect 231646 484718 231882 484954
rect 231326 484398 231562 484634
rect 231646 484398 231882 484634
rect 231326 448718 231562 448954
rect 231646 448718 231882 448954
rect 231326 448398 231562 448634
rect 231646 448398 231882 448634
rect 231326 412718 231562 412954
rect 231646 412718 231882 412954
rect 231326 412398 231562 412634
rect 231646 412398 231882 412634
rect 235826 708442 236062 708678
rect 236146 708442 236382 708678
rect 235826 708122 236062 708358
rect 236146 708122 236382 708358
rect 235826 669218 236062 669454
rect 236146 669218 236382 669454
rect 235826 668898 236062 669134
rect 236146 668898 236382 669134
rect 235826 633218 236062 633454
rect 236146 633218 236382 633454
rect 235826 632898 236062 633134
rect 236146 632898 236382 633134
rect 235826 597218 236062 597454
rect 236146 597218 236382 597454
rect 235826 596898 236062 597134
rect 236146 596898 236382 597134
rect 235826 561218 236062 561454
rect 236146 561218 236382 561454
rect 235826 560898 236062 561134
rect 236146 560898 236382 561134
rect 235826 525218 236062 525454
rect 236146 525218 236382 525454
rect 235826 524898 236062 525134
rect 236146 524898 236382 525134
rect 235826 489218 236062 489454
rect 236146 489218 236382 489454
rect 235826 488898 236062 489134
rect 236146 488898 236382 489134
rect 235826 453218 236062 453454
rect 236146 453218 236382 453454
rect 235826 452898 236062 453134
rect 236146 452898 236382 453134
rect 235826 417218 236062 417454
rect 236146 417218 236382 417454
rect 235826 416898 236062 417134
rect 236146 416898 236382 417134
rect 231326 376718 231562 376954
rect 231646 376718 231882 376954
rect 231326 376398 231562 376634
rect 231646 376398 231882 376634
rect 231326 340718 231562 340954
rect 231646 340718 231882 340954
rect 231326 340398 231562 340634
rect 231646 340398 231882 340634
rect 231326 304718 231562 304954
rect 231646 304718 231882 304954
rect 231326 304398 231562 304634
rect 231646 304398 231882 304634
rect 231326 268718 231562 268954
rect 231646 268718 231882 268954
rect 231326 268398 231562 268634
rect 231646 268398 231882 268634
rect 231326 232718 231562 232954
rect 231646 232718 231882 232954
rect 231326 232398 231562 232634
rect 231646 232398 231882 232634
rect 231326 196718 231562 196954
rect 231646 196718 231882 196954
rect 231326 196398 231562 196634
rect 231646 196398 231882 196634
rect 231326 160718 231562 160954
rect 231646 160718 231882 160954
rect 231326 160398 231562 160634
rect 231646 160398 231882 160634
rect 231326 124718 231562 124954
rect 231646 124718 231882 124954
rect 231326 124398 231562 124634
rect 231646 124398 231882 124634
rect 240326 709402 240562 709638
rect 240646 709402 240882 709638
rect 240326 709082 240562 709318
rect 240646 709082 240882 709318
rect 240326 673718 240562 673954
rect 240646 673718 240882 673954
rect 240326 673398 240562 673634
rect 240646 673398 240882 673634
rect 240326 637718 240562 637954
rect 240646 637718 240882 637954
rect 240326 637398 240562 637634
rect 240646 637398 240882 637634
rect 240326 601718 240562 601954
rect 240646 601718 240882 601954
rect 240326 601398 240562 601634
rect 240646 601398 240882 601634
rect 240326 565718 240562 565954
rect 240646 565718 240882 565954
rect 240326 565398 240562 565634
rect 240646 565398 240882 565634
rect 240326 529718 240562 529954
rect 240646 529718 240882 529954
rect 240326 529398 240562 529634
rect 240646 529398 240882 529634
rect 240326 493718 240562 493954
rect 240646 493718 240882 493954
rect 240326 493398 240562 493634
rect 240646 493398 240882 493634
rect 240326 457718 240562 457954
rect 240646 457718 240882 457954
rect 240326 457398 240562 457634
rect 240646 457398 240882 457634
rect 240326 421718 240562 421954
rect 240646 421718 240882 421954
rect 240326 421398 240562 421634
rect 240646 421398 240882 421634
rect 240326 385718 240562 385954
rect 240646 385718 240882 385954
rect 240326 385398 240562 385634
rect 240646 385398 240882 385634
rect 235826 309218 236062 309454
rect 236146 309218 236382 309454
rect 235826 308898 236062 309134
rect 236146 308898 236382 309134
rect 235826 273218 236062 273454
rect 236146 273218 236382 273454
rect 235826 272898 236062 273134
rect 236146 272898 236382 273134
rect 235826 237218 236062 237454
rect 236146 237218 236382 237454
rect 235826 236898 236062 237134
rect 236146 236898 236382 237134
rect 235826 201218 236062 201454
rect 236146 201218 236382 201454
rect 235826 200898 236062 201134
rect 236146 200898 236382 201134
rect 235826 165218 236062 165454
rect 236146 165218 236382 165454
rect 235826 164898 236062 165134
rect 236146 164898 236382 165134
rect 235826 129218 236062 129454
rect 236146 129218 236382 129454
rect 235826 128898 236062 129134
rect 236146 128898 236382 129134
rect 231326 88718 231562 88954
rect 231646 88718 231882 88954
rect 231326 88398 231562 88634
rect 231646 88398 231882 88634
rect 231326 52718 231562 52954
rect 231646 52718 231882 52954
rect 231326 52398 231562 52634
rect 231646 52398 231882 52634
rect 231326 16718 231562 16954
rect 231646 16718 231882 16954
rect 231326 16398 231562 16634
rect 231646 16398 231882 16634
rect 231326 -3462 231562 -3226
rect 231646 -3462 231882 -3226
rect 231326 -3782 231562 -3546
rect 231646 -3782 231882 -3546
rect 239250 363218 239486 363454
rect 239250 362898 239486 363134
rect 244826 710362 245062 710598
rect 245146 710362 245382 710598
rect 244826 710042 245062 710278
rect 245146 710042 245382 710278
rect 244826 678218 245062 678454
rect 245146 678218 245382 678454
rect 244826 677898 245062 678134
rect 245146 677898 245382 678134
rect 244826 642218 245062 642454
rect 245146 642218 245382 642454
rect 244826 641898 245062 642134
rect 245146 641898 245382 642134
rect 244826 606218 245062 606454
rect 245146 606218 245382 606454
rect 244826 605898 245062 606134
rect 245146 605898 245382 606134
rect 244826 570218 245062 570454
rect 245146 570218 245382 570454
rect 244826 569898 245062 570134
rect 245146 569898 245382 570134
rect 244826 534218 245062 534454
rect 245146 534218 245382 534454
rect 244826 533898 245062 534134
rect 245146 533898 245382 534134
rect 244826 498218 245062 498454
rect 245146 498218 245382 498454
rect 244826 497898 245062 498134
rect 245146 497898 245382 498134
rect 244826 462218 245062 462454
rect 245146 462218 245382 462454
rect 244826 461898 245062 462134
rect 245146 461898 245382 462134
rect 244826 426218 245062 426454
rect 245146 426218 245382 426454
rect 244826 425898 245062 426134
rect 245146 425898 245382 426134
rect 244826 390218 245062 390454
rect 245146 390218 245382 390454
rect 244826 389898 245062 390134
rect 245146 389898 245382 390134
rect 249326 711322 249562 711558
rect 249646 711322 249882 711558
rect 249326 711002 249562 711238
rect 249646 711002 249882 711238
rect 249326 682718 249562 682954
rect 249646 682718 249882 682954
rect 249326 682398 249562 682634
rect 249646 682398 249882 682634
rect 249326 646718 249562 646954
rect 249646 646718 249882 646954
rect 249326 646398 249562 646634
rect 249646 646398 249882 646634
rect 249326 610718 249562 610954
rect 249646 610718 249882 610954
rect 249326 610398 249562 610634
rect 249646 610398 249882 610634
rect 249326 574718 249562 574954
rect 249646 574718 249882 574954
rect 249326 574398 249562 574634
rect 249646 574398 249882 574634
rect 249326 538718 249562 538954
rect 249646 538718 249882 538954
rect 249326 538398 249562 538634
rect 249646 538398 249882 538634
rect 249326 502718 249562 502954
rect 249646 502718 249882 502954
rect 249326 502398 249562 502634
rect 249646 502398 249882 502634
rect 249326 466718 249562 466954
rect 249646 466718 249882 466954
rect 249326 466398 249562 466634
rect 249646 466398 249882 466634
rect 249326 430718 249562 430954
rect 249646 430718 249882 430954
rect 249326 430398 249562 430634
rect 249646 430398 249882 430634
rect 249326 394718 249562 394954
rect 249646 394718 249882 394954
rect 249326 394398 249562 394634
rect 249646 394398 249882 394634
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 253826 651218 254062 651454
rect 254146 651218 254382 651454
rect 253826 650898 254062 651134
rect 254146 650898 254382 651134
rect 253826 615218 254062 615454
rect 254146 615218 254382 615454
rect 253826 614898 254062 615134
rect 254146 614898 254382 615134
rect 253826 579218 254062 579454
rect 254146 579218 254382 579454
rect 253826 578898 254062 579134
rect 254146 578898 254382 579134
rect 253826 543218 254062 543454
rect 254146 543218 254382 543454
rect 253826 542898 254062 543134
rect 254146 542898 254382 543134
rect 253826 507218 254062 507454
rect 254146 507218 254382 507454
rect 253826 506898 254062 507134
rect 254146 506898 254382 507134
rect 253826 471218 254062 471454
rect 254146 471218 254382 471454
rect 253826 470898 254062 471134
rect 254146 470898 254382 471134
rect 253826 435218 254062 435454
rect 254146 435218 254382 435454
rect 253826 434898 254062 435134
rect 254146 434898 254382 435134
rect 253826 399218 254062 399454
rect 254146 399218 254382 399454
rect 253826 398898 254062 399134
rect 254146 398898 254382 399134
rect 258326 705562 258562 705798
rect 258646 705562 258882 705798
rect 258326 705242 258562 705478
rect 258646 705242 258882 705478
rect 258326 691718 258562 691954
rect 258646 691718 258882 691954
rect 258326 691398 258562 691634
rect 258646 691398 258882 691634
rect 258326 655718 258562 655954
rect 258646 655718 258882 655954
rect 258326 655398 258562 655634
rect 258646 655398 258882 655634
rect 258326 619718 258562 619954
rect 258646 619718 258882 619954
rect 258326 619398 258562 619634
rect 258646 619398 258882 619634
rect 258326 583718 258562 583954
rect 258646 583718 258882 583954
rect 258326 583398 258562 583634
rect 258646 583398 258882 583634
rect 258326 547718 258562 547954
rect 258646 547718 258882 547954
rect 258326 547398 258562 547634
rect 258646 547398 258882 547634
rect 258326 511718 258562 511954
rect 258646 511718 258882 511954
rect 258326 511398 258562 511634
rect 258646 511398 258882 511634
rect 258326 475718 258562 475954
rect 258646 475718 258882 475954
rect 258326 475398 258562 475634
rect 258646 475398 258882 475634
rect 258326 439718 258562 439954
rect 258646 439718 258882 439954
rect 258326 439398 258562 439634
rect 258646 439398 258882 439634
rect 258326 403718 258562 403954
rect 258646 403718 258882 403954
rect 258326 403398 258562 403634
rect 258646 403398 258882 403634
rect 262826 706522 263062 706758
rect 263146 706522 263382 706758
rect 262826 706202 263062 706438
rect 263146 706202 263382 706438
rect 262826 696218 263062 696454
rect 263146 696218 263382 696454
rect 262826 695898 263062 696134
rect 263146 695898 263382 696134
rect 262826 660218 263062 660454
rect 263146 660218 263382 660454
rect 262826 659898 263062 660134
rect 263146 659898 263382 660134
rect 262826 624218 263062 624454
rect 263146 624218 263382 624454
rect 262826 623898 263062 624134
rect 263146 623898 263382 624134
rect 262826 588218 263062 588454
rect 263146 588218 263382 588454
rect 262826 587898 263062 588134
rect 263146 587898 263382 588134
rect 262826 552218 263062 552454
rect 263146 552218 263382 552454
rect 262826 551898 263062 552134
rect 263146 551898 263382 552134
rect 262826 516218 263062 516454
rect 263146 516218 263382 516454
rect 262826 515898 263062 516134
rect 263146 515898 263382 516134
rect 262826 480218 263062 480454
rect 263146 480218 263382 480454
rect 262826 479898 263062 480134
rect 263146 479898 263382 480134
rect 262826 444218 263062 444454
rect 263146 444218 263382 444454
rect 262826 443898 263062 444134
rect 263146 443898 263382 444134
rect 262826 408218 263062 408454
rect 263146 408218 263382 408454
rect 262826 407898 263062 408134
rect 263146 407898 263382 408134
rect 267326 707482 267562 707718
rect 267646 707482 267882 707718
rect 267326 707162 267562 707398
rect 267646 707162 267882 707398
rect 267326 700718 267562 700954
rect 267646 700718 267882 700954
rect 267326 700398 267562 700634
rect 267646 700398 267882 700634
rect 267326 664718 267562 664954
rect 267646 664718 267882 664954
rect 267326 664398 267562 664634
rect 267646 664398 267882 664634
rect 267326 628718 267562 628954
rect 267646 628718 267882 628954
rect 267326 628398 267562 628634
rect 267646 628398 267882 628634
rect 267326 592718 267562 592954
rect 267646 592718 267882 592954
rect 267326 592398 267562 592634
rect 267646 592398 267882 592634
rect 267326 556718 267562 556954
rect 267646 556718 267882 556954
rect 267326 556398 267562 556634
rect 267646 556398 267882 556634
rect 267326 520718 267562 520954
rect 267646 520718 267882 520954
rect 267326 520398 267562 520634
rect 267646 520398 267882 520634
rect 267326 484718 267562 484954
rect 267646 484718 267882 484954
rect 267326 484398 267562 484634
rect 267646 484398 267882 484634
rect 267326 448718 267562 448954
rect 267646 448718 267882 448954
rect 267326 448398 267562 448634
rect 267646 448398 267882 448634
rect 267326 412718 267562 412954
rect 267646 412718 267882 412954
rect 267326 412398 267562 412634
rect 267646 412398 267882 412634
rect 271826 708442 272062 708678
rect 272146 708442 272382 708678
rect 271826 708122 272062 708358
rect 272146 708122 272382 708358
rect 271826 669218 272062 669454
rect 272146 669218 272382 669454
rect 271826 668898 272062 669134
rect 272146 668898 272382 669134
rect 271826 633218 272062 633454
rect 272146 633218 272382 633454
rect 271826 632898 272062 633134
rect 272146 632898 272382 633134
rect 271826 597218 272062 597454
rect 272146 597218 272382 597454
rect 271826 596898 272062 597134
rect 272146 596898 272382 597134
rect 271826 561218 272062 561454
rect 272146 561218 272382 561454
rect 271826 560898 272062 561134
rect 272146 560898 272382 561134
rect 271826 525218 272062 525454
rect 272146 525218 272382 525454
rect 271826 524898 272062 525134
rect 272146 524898 272382 525134
rect 271826 489218 272062 489454
rect 272146 489218 272382 489454
rect 271826 488898 272062 489134
rect 272146 488898 272382 489134
rect 271826 453218 272062 453454
rect 272146 453218 272382 453454
rect 271826 452898 272062 453134
rect 272146 452898 272382 453134
rect 271826 417218 272062 417454
rect 272146 417218 272382 417454
rect 271826 416898 272062 417134
rect 272146 416898 272382 417134
rect 276326 709402 276562 709638
rect 276646 709402 276882 709638
rect 276326 709082 276562 709318
rect 276646 709082 276882 709318
rect 276326 673718 276562 673954
rect 276646 673718 276882 673954
rect 276326 673398 276562 673634
rect 276646 673398 276882 673634
rect 276326 637718 276562 637954
rect 276646 637718 276882 637954
rect 276326 637398 276562 637634
rect 276646 637398 276882 637634
rect 276326 601718 276562 601954
rect 276646 601718 276882 601954
rect 276326 601398 276562 601634
rect 276646 601398 276882 601634
rect 276326 565718 276562 565954
rect 276646 565718 276882 565954
rect 276326 565398 276562 565634
rect 276646 565398 276882 565634
rect 276326 529718 276562 529954
rect 276646 529718 276882 529954
rect 276326 529398 276562 529634
rect 276646 529398 276882 529634
rect 276326 493718 276562 493954
rect 276646 493718 276882 493954
rect 276326 493398 276562 493634
rect 276646 493398 276882 493634
rect 276326 457718 276562 457954
rect 276646 457718 276882 457954
rect 276326 457398 276562 457634
rect 276646 457398 276882 457634
rect 276326 421718 276562 421954
rect 276646 421718 276882 421954
rect 276326 421398 276562 421634
rect 276646 421398 276882 421634
rect 276326 385718 276562 385954
rect 276646 385718 276882 385954
rect 276326 385398 276562 385634
rect 276646 385398 276882 385634
rect 280826 710362 281062 710598
rect 281146 710362 281382 710598
rect 280826 710042 281062 710278
rect 281146 710042 281382 710278
rect 280826 678218 281062 678454
rect 281146 678218 281382 678454
rect 280826 677898 281062 678134
rect 281146 677898 281382 678134
rect 280826 642218 281062 642454
rect 281146 642218 281382 642454
rect 280826 641898 281062 642134
rect 281146 641898 281382 642134
rect 280826 606218 281062 606454
rect 281146 606218 281382 606454
rect 280826 605898 281062 606134
rect 281146 605898 281382 606134
rect 280826 570218 281062 570454
rect 281146 570218 281382 570454
rect 280826 569898 281062 570134
rect 281146 569898 281382 570134
rect 280826 534218 281062 534454
rect 281146 534218 281382 534454
rect 280826 533898 281062 534134
rect 281146 533898 281382 534134
rect 280826 498218 281062 498454
rect 281146 498218 281382 498454
rect 280826 497898 281062 498134
rect 281146 497898 281382 498134
rect 280826 462218 281062 462454
rect 281146 462218 281382 462454
rect 280826 461898 281062 462134
rect 281146 461898 281382 462134
rect 280826 426218 281062 426454
rect 281146 426218 281382 426454
rect 280826 425898 281062 426134
rect 281146 425898 281382 426134
rect 280826 390218 281062 390454
rect 281146 390218 281382 390454
rect 280826 389898 281062 390134
rect 281146 389898 281382 390134
rect 285326 711322 285562 711558
rect 285646 711322 285882 711558
rect 285326 711002 285562 711238
rect 285646 711002 285882 711238
rect 285326 682718 285562 682954
rect 285646 682718 285882 682954
rect 285326 682398 285562 682634
rect 285646 682398 285882 682634
rect 285326 646718 285562 646954
rect 285646 646718 285882 646954
rect 285326 646398 285562 646634
rect 285646 646398 285882 646634
rect 285326 610718 285562 610954
rect 285646 610718 285882 610954
rect 285326 610398 285562 610634
rect 285646 610398 285882 610634
rect 285326 574718 285562 574954
rect 285646 574718 285882 574954
rect 285326 574398 285562 574634
rect 285646 574398 285882 574634
rect 285326 538718 285562 538954
rect 285646 538718 285882 538954
rect 285326 538398 285562 538634
rect 285646 538398 285882 538634
rect 285326 502718 285562 502954
rect 285646 502718 285882 502954
rect 285326 502398 285562 502634
rect 285646 502398 285882 502634
rect 285326 466718 285562 466954
rect 285646 466718 285882 466954
rect 285326 466398 285562 466634
rect 285646 466398 285882 466634
rect 285326 430718 285562 430954
rect 285646 430718 285882 430954
rect 285326 430398 285562 430634
rect 285646 430398 285882 430634
rect 285326 394718 285562 394954
rect 285646 394718 285882 394954
rect 285326 394398 285562 394634
rect 285646 394398 285882 394634
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 289826 651218 290062 651454
rect 290146 651218 290382 651454
rect 289826 650898 290062 651134
rect 290146 650898 290382 651134
rect 289826 615218 290062 615454
rect 290146 615218 290382 615454
rect 289826 614898 290062 615134
rect 290146 614898 290382 615134
rect 289826 579218 290062 579454
rect 290146 579218 290382 579454
rect 289826 578898 290062 579134
rect 290146 578898 290382 579134
rect 289826 543218 290062 543454
rect 290146 543218 290382 543454
rect 289826 542898 290062 543134
rect 290146 542898 290382 543134
rect 289826 507218 290062 507454
rect 290146 507218 290382 507454
rect 289826 506898 290062 507134
rect 290146 506898 290382 507134
rect 289826 471218 290062 471454
rect 290146 471218 290382 471454
rect 289826 470898 290062 471134
rect 290146 470898 290382 471134
rect 289826 435218 290062 435454
rect 290146 435218 290382 435454
rect 289826 434898 290062 435134
rect 290146 434898 290382 435134
rect 289826 399218 290062 399454
rect 290146 399218 290382 399454
rect 289826 398898 290062 399134
rect 290146 398898 290382 399134
rect 294326 705562 294562 705798
rect 294646 705562 294882 705798
rect 294326 705242 294562 705478
rect 294646 705242 294882 705478
rect 294326 691718 294562 691954
rect 294646 691718 294882 691954
rect 294326 691398 294562 691634
rect 294646 691398 294882 691634
rect 294326 655718 294562 655954
rect 294646 655718 294882 655954
rect 294326 655398 294562 655634
rect 294646 655398 294882 655634
rect 294326 619718 294562 619954
rect 294646 619718 294882 619954
rect 294326 619398 294562 619634
rect 294646 619398 294882 619634
rect 294326 583718 294562 583954
rect 294646 583718 294882 583954
rect 294326 583398 294562 583634
rect 294646 583398 294882 583634
rect 294326 547718 294562 547954
rect 294646 547718 294882 547954
rect 294326 547398 294562 547634
rect 294646 547398 294882 547634
rect 294326 511718 294562 511954
rect 294646 511718 294882 511954
rect 294326 511398 294562 511634
rect 294646 511398 294882 511634
rect 294326 475718 294562 475954
rect 294646 475718 294882 475954
rect 294326 475398 294562 475634
rect 294646 475398 294882 475634
rect 294326 439718 294562 439954
rect 294646 439718 294882 439954
rect 294326 439398 294562 439634
rect 294646 439398 294882 439634
rect 294326 403718 294562 403954
rect 294646 403718 294882 403954
rect 294326 403398 294562 403634
rect 294646 403398 294882 403634
rect 254610 367718 254846 367954
rect 254610 367398 254846 367634
rect 285330 367718 285566 367954
rect 285330 367398 285566 367634
rect 269970 363218 270206 363454
rect 269970 362898 270206 363134
rect 240326 313718 240562 313954
rect 240646 313718 240882 313954
rect 240326 313398 240562 313634
rect 240646 313398 240882 313634
rect 240326 277718 240562 277954
rect 240646 277718 240882 277954
rect 240326 277398 240562 277634
rect 240646 277398 240882 277634
rect 240326 241718 240562 241954
rect 240646 241718 240882 241954
rect 240326 241398 240562 241634
rect 240646 241398 240882 241634
rect 240326 205718 240562 205954
rect 240646 205718 240882 205954
rect 240326 205398 240562 205634
rect 240646 205398 240882 205634
rect 240326 169718 240562 169954
rect 240646 169718 240882 169954
rect 240326 169398 240562 169634
rect 240646 169398 240882 169634
rect 240326 133718 240562 133954
rect 240646 133718 240882 133954
rect 240326 133398 240562 133634
rect 240646 133398 240882 133634
rect 240326 97718 240562 97954
rect 240646 97718 240882 97954
rect 235826 93218 236062 93454
rect 236146 93218 236382 93454
rect 235826 92898 236062 93134
rect 236146 92898 236382 93134
rect 235826 57218 236062 57454
rect 236146 57218 236382 57454
rect 235826 56898 236062 57134
rect 236146 56898 236382 57134
rect 235826 21218 236062 21454
rect 236146 21218 236382 21454
rect 235826 20898 236062 21134
rect 236146 20898 236382 21134
rect 235826 -4422 236062 -4186
rect 236146 -4422 236382 -4186
rect 235826 -4742 236062 -4506
rect 236146 -4742 236382 -4506
rect 240326 97398 240562 97634
rect 240646 97398 240882 97634
rect 240326 61718 240562 61954
rect 240646 61718 240882 61954
rect 240326 61398 240562 61634
rect 240646 61398 240882 61634
rect 240326 25718 240562 25954
rect 240646 25718 240882 25954
rect 240326 25398 240562 25634
rect 240646 25398 240882 25634
rect 244826 318218 245062 318454
rect 245146 318218 245382 318454
rect 244826 317898 245062 318134
rect 245146 317898 245382 318134
rect 244826 282218 245062 282454
rect 245146 282218 245382 282454
rect 244826 281898 245062 282134
rect 245146 281898 245382 282134
rect 244826 246218 245062 246454
rect 245146 246218 245382 246454
rect 244826 245898 245062 246134
rect 245146 245898 245382 246134
rect 244826 210218 245062 210454
rect 245146 210218 245382 210454
rect 244826 209898 245062 210134
rect 245146 209898 245382 210134
rect 244826 174218 245062 174454
rect 245146 174218 245382 174454
rect 244826 173898 245062 174134
rect 245146 173898 245382 174134
rect 244826 138218 245062 138454
rect 245146 138218 245382 138454
rect 244826 137898 245062 138134
rect 245146 137898 245382 138134
rect 244826 102218 245062 102454
rect 245146 102218 245382 102454
rect 244826 101898 245062 102134
rect 245146 101898 245382 102134
rect 244826 66218 245062 66454
rect 245146 66218 245382 66454
rect 244826 65898 245062 66134
rect 245146 65898 245382 66134
rect 244826 30218 245062 30454
rect 245146 30218 245382 30454
rect 244826 29898 245062 30134
rect 245146 29898 245382 30134
rect 240326 -5382 240562 -5146
rect 240646 -5382 240882 -5146
rect 240326 -5702 240562 -5466
rect 240646 -5702 240882 -5466
rect 249326 322718 249562 322954
rect 249646 322718 249882 322954
rect 249326 322398 249562 322634
rect 249646 322398 249882 322634
rect 249326 286718 249562 286954
rect 249646 286718 249882 286954
rect 249326 286398 249562 286634
rect 249646 286398 249882 286634
rect 249326 250718 249562 250954
rect 249646 250718 249882 250954
rect 249326 250398 249562 250634
rect 249646 250398 249882 250634
rect 249326 214718 249562 214954
rect 249646 214718 249882 214954
rect 249326 214398 249562 214634
rect 249646 214398 249882 214634
rect 249326 178718 249562 178954
rect 249646 178718 249882 178954
rect 249326 178398 249562 178634
rect 249646 178398 249882 178634
rect 249326 142718 249562 142954
rect 249646 142718 249882 142954
rect 249326 142398 249562 142634
rect 249646 142398 249882 142634
rect 249326 106718 249562 106954
rect 249646 106718 249882 106954
rect 249326 106398 249562 106634
rect 249646 106398 249882 106634
rect 249326 70718 249562 70954
rect 249646 70718 249882 70954
rect 249326 70398 249562 70634
rect 249646 70398 249882 70634
rect 249326 34718 249562 34954
rect 249646 34718 249882 34954
rect 249326 34398 249562 34634
rect 249646 34398 249882 34634
rect 244826 -6342 245062 -6106
rect 245146 -6342 245382 -6106
rect 244826 -6662 245062 -6426
rect 245146 -6662 245382 -6426
rect 253826 327218 254062 327454
rect 254146 327218 254382 327454
rect 253826 326898 254062 327134
rect 254146 326898 254382 327134
rect 253826 291218 254062 291454
rect 254146 291218 254382 291454
rect 253826 290898 254062 291134
rect 254146 290898 254382 291134
rect 253826 255218 254062 255454
rect 254146 255218 254382 255454
rect 253826 254898 254062 255134
rect 254146 254898 254382 255134
rect 253826 219218 254062 219454
rect 254146 219218 254382 219454
rect 253826 218898 254062 219134
rect 254146 218898 254382 219134
rect 253826 183218 254062 183454
rect 254146 183218 254382 183454
rect 253826 182898 254062 183134
rect 254146 182898 254382 183134
rect 253826 147218 254062 147454
rect 254146 147218 254382 147454
rect 253826 146898 254062 147134
rect 254146 146898 254382 147134
rect 253826 111218 254062 111454
rect 254146 111218 254382 111454
rect 253826 110898 254062 111134
rect 254146 110898 254382 111134
rect 253826 75218 254062 75454
rect 254146 75218 254382 75454
rect 253826 74898 254062 75134
rect 254146 74898 254382 75134
rect 253826 39218 254062 39454
rect 254146 39218 254382 39454
rect 253826 38898 254062 39134
rect 254146 38898 254382 39134
rect 249326 -7302 249562 -7066
rect 249646 -7302 249882 -7066
rect 249326 -7622 249562 -7386
rect 249646 -7622 249882 -7386
rect 258326 331718 258562 331954
rect 258646 331718 258882 331954
rect 258326 331398 258562 331634
rect 258646 331398 258882 331634
rect 258326 295718 258562 295954
rect 258646 295718 258882 295954
rect 258326 295398 258562 295634
rect 258646 295398 258882 295634
rect 258326 259718 258562 259954
rect 258646 259718 258882 259954
rect 258326 259398 258562 259634
rect 258646 259398 258882 259634
rect 258326 223718 258562 223954
rect 258646 223718 258882 223954
rect 258326 223398 258562 223634
rect 258646 223398 258882 223634
rect 258326 187718 258562 187954
rect 258646 187718 258882 187954
rect 258326 187398 258562 187634
rect 258646 187398 258882 187634
rect 258326 79718 258562 79954
rect 258646 79718 258882 79954
rect 258326 79398 258562 79634
rect 258646 79398 258882 79634
rect 258326 43718 258562 43954
rect 258646 43718 258882 43954
rect 258326 43398 258562 43634
rect 258646 43398 258882 43634
rect 258326 7718 258562 7954
rect 258646 7718 258882 7954
rect 258326 7398 258562 7634
rect 258646 7398 258882 7634
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 262826 300218 263062 300454
rect 263146 300218 263382 300454
rect 262826 299898 263062 300134
rect 263146 299898 263382 300134
rect 262826 264218 263062 264454
rect 263146 264218 263382 264454
rect 262826 263898 263062 264134
rect 263146 263898 263382 264134
rect 262826 228218 263062 228454
rect 263146 228218 263382 228454
rect 262826 227898 263062 228134
rect 263146 227898 263382 228134
rect 262826 192218 263062 192454
rect 263146 192218 263382 192454
rect 262826 191898 263062 192134
rect 263146 191898 263382 192134
rect 267326 304718 267562 304954
rect 267646 304718 267882 304954
rect 267326 304398 267562 304634
rect 267646 304398 267882 304634
rect 267326 268718 267562 268954
rect 267646 268718 267882 268954
rect 267326 268398 267562 268634
rect 267646 268398 267882 268634
rect 267326 232718 267562 232954
rect 267646 232718 267882 232954
rect 267326 232398 267562 232634
rect 267646 232398 267882 232634
rect 267326 196718 267562 196954
rect 267646 196718 267882 196954
rect 267326 196398 267562 196634
rect 267646 196398 267882 196634
rect 267326 160718 267562 160954
rect 267646 160718 267882 160954
rect 267326 160398 267562 160634
rect 267646 160398 267882 160634
rect 271826 309218 272062 309454
rect 272146 309218 272382 309454
rect 271826 308898 272062 309134
rect 272146 308898 272382 309134
rect 271826 273218 272062 273454
rect 272146 273218 272382 273454
rect 271826 272898 272062 273134
rect 272146 272898 272382 273134
rect 271826 237218 272062 237454
rect 272146 237218 272382 237454
rect 271826 236898 272062 237134
rect 272146 236898 272382 237134
rect 271826 201218 272062 201454
rect 272146 201218 272382 201454
rect 271826 200898 272062 201134
rect 272146 200898 272382 201134
rect 271826 165218 272062 165454
rect 272146 165218 272382 165454
rect 271826 164898 272062 165134
rect 272146 164898 272382 165134
rect 276326 313718 276562 313954
rect 276646 313718 276882 313954
rect 276326 313398 276562 313634
rect 276646 313398 276882 313634
rect 276326 277718 276562 277954
rect 276646 277718 276882 277954
rect 276326 277398 276562 277634
rect 276646 277398 276882 277634
rect 276326 241718 276562 241954
rect 276646 241718 276882 241954
rect 276326 241398 276562 241634
rect 276646 241398 276882 241634
rect 276326 205718 276562 205954
rect 276646 205718 276882 205954
rect 276326 205398 276562 205634
rect 276646 205398 276882 205634
rect 276326 169718 276562 169954
rect 276646 169718 276882 169954
rect 276326 169398 276562 169634
rect 276646 169398 276882 169634
rect 280826 318218 281062 318454
rect 281146 318218 281382 318454
rect 280826 317898 281062 318134
rect 281146 317898 281382 318134
rect 280826 282218 281062 282454
rect 281146 282218 281382 282454
rect 280826 281898 281062 282134
rect 281146 281898 281382 282134
rect 280826 246218 281062 246454
rect 281146 246218 281382 246454
rect 280826 245898 281062 246134
rect 281146 245898 281382 246134
rect 280826 210218 281062 210454
rect 281146 210218 281382 210454
rect 280826 209898 281062 210134
rect 281146 209898 281382 210134
rect 280826 174218 281062 174454
rect 281146 174218 281382 174454
rect 280826 173898 281062 174134
rect 281146 173898 281382 174134
rect 285326 322718 285562 322954
rect 285646 322718 285882 322954
rect 285326 322398 285562 322634
rect 285646 322398 285882 322634
rect 285326 286718 285562 286954
rect 285646 286718 285882 286954
rect 285326 286398 285562 286634
rect 285646 286398 285882 286634
rect 285326 250718 285562 250954
rect 285646 250718 285882 250954
rect 285326 250398 285562 250634
rect 285646 250398 285882 250634
rect 285326 214718 285562 214954
rect 285646 214718 285882 214954
rect 285326 214398 285562 214634
rect 285646 214398 285882 214634
rect 285326 178718 285562 178954
rect 285646 178718 285882 178954
rect 285326 178398 285562 178634
rect 285646 178398 285882 178634
rect 289826 327218 290062 327454
rect 290146 327218 290382 327454
rect 289826 326898 290062 327134
rect 290146 326898 290382 327134
rect 289826 291218 290062 291454
rect 290146 291218 290382 291454
rect 289826 290898 290062 291134
rect 290146 290898 290382 291134
rect 289826 255218 290062 255454
rect 290146 255218 290382 255454
rect 289826 254898 290062 255134
rect 290146 254898 290382 255134
rect 289826 219218 290062 219454
rect 290146 219218 290382 219454
rect 289826 218898 290062 219134
rect 290146 218898 290382 219134
rect 289826 183218 290062 183454
rect 290146 183218 290382 183454
rect 289826 182898 290062 183134
rect 290146 182898 290382 183134
rect 298826 706522 299062 706758
rect 299146 706522 299382 706758
rect 298826 706202 299062 706438
rect 299146 706202 299382 706438
rect 298826 696218 299062 696454
rect 299146 696218 299382 696454
rect 298826 695898 299062 696134
rect 299146 695898 299382 696134
rect 298826 660218 299062 660454
rect 299146 660218 299382 660454
rect 298826 659898 299062 660134
rect 299146 659898 299382 660134
rect 298826 624218 299062 624454
rect 299146 624218 299382 624454
rect 298826 623898 299062 624134
rect 299146 623898 299382 624134
rect 298826 588218 299062 588454
rect 299146 588218 299382 588454
rect 298826 587898 299062 588134
rect 299146 587898 299382 588134
rect 298826 552218 299062 552454
rect 299146 552218 299382 552454
rect 298826 551898 299062 552134
rect 299146 551898 299382 552134
rect 298826 516218 299062 516454
rect 299146 516218 299382 516454
rect 298826 515898 299062 516134
rect 299146 515898 299382 516134
rect 298826 480218 299062 480454
rect 299146 480218 299382 480454
rect 298826 479898 299062 480134
rect 299146 479898 299382 480134
rect 298826 444218 299062 444454
rect 299146 444218 299382 444454
rect 298826 443898 299062 444134
rect 299146 443898 299382 444134
rect 298826 408218 299062 408454
rect 299146 408218 299382 408454
rect 298826 407898 299062 408134
rect 299146 407898 299382 408134
rect 294326 331718 294562 331954
rect 294646 331718 294882 331954
rect 294326 331398 294562 331634
rect 294646 331398 294882 331634
rect 294326 295718 294562 295954
rect 294646 295718 294882 295954
rect 294326 295398 294562 295634
rect 294646 295398 294882 295634
rect 294326 259718 294562 259954
rect 294646 259718 294882 259954
rect 294326 259398 294562 259634
rect 294646 259398 294882 259634
rect 294326 223718 294562 223954
rect 294646 223718 294882 223954
rect 294326 223398 294562 223634
rect 294646 223398 294882 223634
rect 294326 187718 294562 187954
rect 294646 187718 294882 187954
rect 294326 187398 294562 187634
rect 294646 187398 294882 187634
rect 303326 707482 303562 707718
rect 303646 707482 303882 707718
rect 303326 707162 303562 707398
rect 303646 707162 303882 707398
rect 303326 700718 303562 700954
rect 303646 700718 303882 700954
rect 303326 700398 303562 700634
rect 303646 700398 303882 700634
rect 303326 664718 303562 664954
rect 303646 664718 303882 664954
rect 303326 664398 303562 664634
rect 303646 664398 303882 664634
rect 303326 628718 303562 628954
rect 303646 628718 303882 628954
rect 303326 628398 303562 628634
rect 303646 628398 303882 628634
rect 303326 592718 303562 592954
rect 303646 592718 303882 592954
rect 303326 592398 303562 592634
rect 303646 592398 303882 592634
rect 303326 556718 303562 556954
rect 303646 556718 303882 556954
rect 303326 556398 303562 556634
rect 303646 556398 303882 556634
rect 303326 520718 303562 520954
rect 303646 520718 303882 520954
rect 303326 520398 303562 520634
rect 303646 520398 303882 520634
rect 303326 484718 303562 484954
rect 303646 484718 303882 484954
rect 303326 484398 303562 484634
rect 303646 484398 303882 484634
rect 303326 448718 303562 448954
rect 303646 448718 303882 448954
rect 303326 448398 303562 448634
rect 303646 448398 303882 448634
rect 303326 412718 303562 412954
rect 303646 412718 303882 412954
rect 303326 412398 303562 412634
rect 303646 412398 303882 412634
rect 303326 376718 303562 376954
rect 303646 376718 303882 376954
rect 303326 376398 303562 376634
rect 303646 376398 303882 376634
rect 303326 340718 303562 340954
rect 303646 340718 303882 340954
rect 303326 340398 303562 340634
rect 303646 340398 303882 340634
rect 298826 300218 299062 300454
rect 299146 300218 299382 300454
rect 298826 299898 299062 300134
rect 299146 299898 299382 300134
rect 298826 264218 299062 264454
rect 299146 264218 299382 264454
rect 298826 263898 299062 264134
rect 299146 263898 299382 264134
rect 298826 228218 299062 228454
rect 299146 228218 299382 228454
rect 298826 227898 299062 228134
rect 299146 227898 299382 228134
rect 298826 192218 299062 192454
rect 299146 192218 299382 192454
rect 298826 191898 299062 192134
rect 299146 191898 299382 192134
rect 303326 304718 303562 304954
rect 303646 304718 303882 304954
rect 303326 304398 303562 304634
rect 303646 304398 303882 304634
rect 303326 268718 303562 268954
rect 303646 268718 303882 268954
rect 303326 268398 303562 268634
rect 303646 268398 303882 268634
rect 303326 232718 303562 232954
rect 303646 232718 303882 232954
rect 303326 232398 303562 232634
rect 303646 232398 303882 232634
rect 303326 196718 303562 196954
rect 303646 196718 303882 196954
rect 303326 196398 303562 196634
rect 303646 196398 303882 196634
rect 303326 160718 303562 160954
rect 303646 160718 303882 160954
rect 303326 160398 303562 160634
rect 303646 160398 303882 160634
rect 307826 708442 308062 708678
rect 308146 708442 308382 708678
rect 307826 708122 308062 708358
rect 308146 708122 308382 708358
rect 307826 669218 308062 669454
rect 308146 669218 308382 669454
rect 307826 668898 308062 669134
rect 308146 668898 308382 669134
rect 307826 633218 308062 633454
rect 308146 633218 308382 633454
rect 307826 632898 308062 633134
rect 308146 632898 308382 633134
rect 307826 597218 308062 597454
rect 308146 597218 308382 597454
rect 307826 596898 308062 597134
rect 308146 596898 308382 597134
rect 307826 561218 308062 561454
rect 308146 561218 308382 561454
rect 307826 560898 308062 561134
rect 308146 560898 308382 561134
rect 307826 525218 308062 525454
rect 308146 525218 308382 525454
rect 307826 524898 308062 525134
rect 308146 524898 308382 525134
rect 307826 489218 308062 489454
rect 308146 489218 308382 489454
rect 307826 488898 308062 489134
rect 308146 488898 308382 489134
rect 307826 453218 308062 453454
rect 308146 453218 308382 453454
rect 307826 452898 308062 453134
rect 308146 452898 308382 453134
rect 307826 417218 308062 417454
rect 308146 417218 308382 417454
rect 307826 416898 308062 417134
rect 308146 416898 308382 417134
rect 307826 381218 308062 381454
rect 308146 381218 308382 381454
rect 307826 380898 308062 381134
rect 308146 380898 308382 381134
rect 307826 345218 308062 345454
rect 308146 345218 308382 345454
rect 307826 344898 308062 345134
rect 308146 344898 308382 345134
rect 307826 309218 308062 309454
rect 308146 309218 308382 309454
rect 307826 308898 308062 309134
rect 308146 308898 308382 309134
rect 307826 273218 308062 273454
rect 308146 273218 308382 273454
rect 307826 272898 308062 273134
rect 308146 272898 308382 273134
rect 307826 237218 308062 237454
rect 308146 237218 308382 237454
rect 307826 236898 308062 237134
rect 308146 236898 308382 237134
rect 307826 201218 308062 201454
rect 308146 201218 308382 201454
rect 307826 200898 308062 201134
rect 308146 200898 308382 201134
rect 307826 165218 308062 165454
rect 308146 165218 308382 165454
rect 307826 164898 308062 165134
rect 308146 164898 308382 165134
rect 312326 709402 312562 709638
rect 312646 709402 312882 709638
rect 312326 709082 312562 709318
rect 312646 709082 312882 709318
rect 312326 673718 312562 673954
rect 312646 673718 312882 673954
rect 312326 673398 312562 673634
rect 312646 673398 312882 673634
rect 312326 637718 312562 637954
rect 312646 637718 312882 637954
rect 312326 637398 312562 637634
rect 312646 637398 312882 637634
rect 312326 601718 312562 601954
rect 312646 601718 312882 601954
rect 312326 601398 312562 601634
rect 312646 601398 312882 601634
rect 312326 565718 312562 565954
rect 312646 565718 312882 565954
rect 312326 565398 312562 565634
rect 312646 565398 312882 565634
rect 312326 529718 312562 529954
rect 312646 529718 312882 529954
rect 312326 529398 312562 529634
rect 312646 529398 312882 529634
rect 312326 493718 312562 493954
rect 312646 493718 312882 493954
rect 312326 493398 312562 493634
rect 312646 493398 312882 493634
rect 312326 457718 312562 457954
rect 312646 457718 312882 457954
rect 312326 457398 312562 457634
rect 312646 457398 312882 457634
rect 312326 421718 312562 421954
rect 312646 421718 312882 421954
rect 312326 421398 312562 421634
rect 312646 421398 312882 421634
rect 312326 385718 312562 385954
rect 312646 385718 312882 385954
rect 312326 385398 312562 385634
rect 312646 385398 312882 385634
rect 312326 349718 312562 349954
rect 312646 349718 312882 349954
rect 312326 349398 312562 349634
rect 312646 349398 312882 349634
rect 312326 313718 312562 313954
rect 312646 313718 312882 313954
rect 312326 313398 312562 313634
rect 312646 313398 312882 313634
rect 312326 277718 312562 277954
rect 312646 277718 312882 277954
rect 312326 277398 312562 277634
rect 312646 277398 312882 277634
rect 312326 241718 312562 241954
rect 312646 241718 312882 241954
rect 312326 241398 312562 241634
rect 312646 241398 312882 241634
rect 312326 205718 312562 205954
rect 312646 205718 312882 205954
rect 312326 205398 312562 205634
rect 312646 205398 312882 205634
rect 312326 169718 312562 169954
rect 312646 169718 312882 169954
rect 312326 169398 312562 169634
rect 312646 169398 312882 169634
rect 316826 710362 317062 710598
rect 317146 710362 317382 710598
rect 316826 710042 317062 710278
rect 317146 710042 317382 710278
rect 316826 678218 317062 678454
rect 317146 678218 317382 678454
rect 316826 677898 317062 678134
rect 317146 677898 317382 678134
rect 316826 642218 317062 642454
rect 317146 642218 317382 642454
rect 316826 641898 317062 642134
rect 317146 641898 317382 642134
rect 316826 606218 317062 606454
rect 317146 606218 317382 606454
rect 316826 605898 317062 606134
rect 317146 605898 317382 606134
rect 316826 570218 317062 570454
rect 317146 570218 317382 570454
rect 316826 569898 317062 570134
rect 317146 569898 317382 570134
rect 316826 534218 317062 534454
rect 317146 534218 317382 534454
rect 316826 533898 317062 534134
rect 317146 533898 317382 534134
rect 316826 498218 317062 498454
rect 317146 498218 317382 498454
rect 316826 497898 317062 498134
rect 317146 497898 317382 498134
rect 316826 462218 317062 462454
rect 317146 462218 317382 462454
rect 316826 461898 317062 462134
rect 317146 461898 317382 462134
rect 316826 426218 317062 426454
rect 317146 426218 317382 426454
rect 316826 425898 317062 426134
rect 317146 425898 317382 426134
rect 316826 390218 317062 390454
rect 317146 390218 317382 390454
rect 316826 389898 317062 390134
rect 317146 389898 317382 390134
rect 316826 354218 317062 354454
rect 317146 354218 317382 354454
rect 316826 353898 317062 354134
rect 317146 353898 317382 354134
rect 316826 318218 317062 318454
rect 317146 318218 317382 318454
rect 316826 317898 317062 318134
rect 317146 317898 317382 318134
rect 316826 282218 317062 282454
rect 317146 282218 317382 282454
rect 316826 281898 317062 282134
rect 317146 281898 317382 282134
rect 316826 246218 317062 246454
rect 317146 246218 317382 246454
rect 316826 245898 317062 246134
rect 317146 245898 317382 246134
rect 316826 210218 317062 210454
rect 317146 210218 317382 210454
rect 316826 209898 317062 210134
rect 317146 209898 317382 210134
rect 316826 174218 317062 174454
rect 317146 174218 317382 174454
rect 316826 173898 317062 174134
rect 317146 173898 317382 174134
rect 321326 711322 321562 711558
rect 321646 711322 321882 711558
rect 321326 711002 321562 711238
rect 321646 711002 321882 711238
rect 321326 682718 321562 682954
rect 321646 682718 321882 682954
rect 321326 682398 321562 682634
rect 321646 682398 321882 682634
rect 321326 646718 321562 646954
rect 321646 646718 321882 646954
rect 321326 646398 321562 646634
rect 321646 646398 321882 646634
rect 321326 610718 321562 610954
rect 321646 610718 321882 610954
rect 321326 610398 321562 610634
rect 321646 610398 321882 610634
rect 321326 574718 321562 574954
rect 321646 574718 321882 574954
rect 321326 574398 321562 574634
rect 321646 574398 321882 574634
rect 321326 538718 321562 538954
rect 321646 538718 321882 538954
rect 321326 538398 321562 538634
rect 321646 538398 321882 538634
rect 321326 502718 321562 502954
rect 321646 502718 321882 502954
rect 321326 502398 321562 502634
rect 321646 502398 321882 502634
rect 321326 466718 321562 466954
rect 321646 466718 321882 466954
rect 321326 466398 321562 466634
rect 321646 466398 321882 466634
rect 321326 430718 321562 430954
rect 321646 430718 321882 430954
rect 321326 430398 321562 430634
rect 321646 430398 321882 430634
rect 321326 394718 321562 394954
rect 321646 394718 321882 394954
rect 321326 394398 321562 394634
rect 321646 394398 321882 394634
rect 321326 358718 321562 358954
rect 321646 358718 321882 358954
rect 321326 358398 321562 358634
rect 321646 358398 321882 358634
rect 321326 322718 321562 322954
rect 321646 322718 321882 322954
rect 321326 322398 321562 322634
rect 321646 322398 321882 322634
rect 321326 286718 321562 286954
rect 321646 286718 321882 286954
rect 321326 286398 321562 286634
rect 321646 286398 321882 286634
rect 321326 250718 321562 250954
rect 321646 250718 321882 250954
rect 321326 250398 321562 250634
rect 321646 250398 321882 250634
rect 321326 214718 321562 214954
rect 321646 214718 321882 214954
rect 321326 214398 321562 214634
rect 321646 214398 321882 214634
rect 321326 178718 321562 178954
rect 321646 178718 321882 178954
rect 321326 178398 321562 178634
rect 321646 178398 321882 178634
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 325826 651218 326062 651454
rect 326146 651218 326382 651454
rect 325826 650898 326062 651134
rect 326146 650898 326382 651134
rect 325826 615218 326062 615454
rect 326146 615218 326382 615454
rect 325826 614898 326062 615134
rect 326146 614898 326382 615134
rect 325826 579218 326062 579454
rect 326146 579218 326382 579454
rect 325826 578898 326062 579134
rect 326146 578898 326382 579134
rect 325826 543218 326062 543454
rect 326146 543218 326382 543454
rect 325826 542898 326062 543134
rect 326146 542898 326382 543134
rect 325826 507218 326062 507454
rect 326146 507218 326382 507454
rect 325826 506898 326062 507134
rect 326146 506898 326382 507134
rect 325826 471218 326062 471454
rect 326146 471218 326382 471454
rect 325826 470898 326062 471134
rect 326146 470898 326382 471134
rect 325826 435218 326062 435454
rect 326146 435218 326382 435454
rect 325826 434898 326062 435134
rect 326146 434898 326382 435134
rect 325826 399218 326062 399454
rect 326146 399218 326382 399454
rect 325826 398898 326062 399134
rect 326146 398898 326382 399134
rect 325826 363218 326062 363454
rect 326146 363218 326382 363454
rect 325826 362898 326062 363134
rect 326146 362898 326382 363134
rect 325826 327218 326062 327454
rect 326146 327218 326382 327454
rect 325826 326898 326062 327134
rect 326146 326898 326382 327134
rect 325826 291218 326062 291454
rect 326146 291218 326382 291454
rect 325826 290898 326062 291134
rect 326146 290898 326382 291134
rect 325826 255218 326062 255454
rect 326146 255218 326382 255454
rect 325826 254898 326062 255134
rect 326146 254898 326382 255134
rect 325826 219218 326062 219454
rect 326146 219218 326382 219454
rect 325826 218898 326062 219134
rect 326146 218898 326382 219134
rect 325826 183218 326062 183454
rect 326146 183218 326382 183454
rect 325826 182898 326062 183134
rect 326146 182898 326382 183134
rect 330326 705562 330562 705798
rect 330646 705562 330882 705798
rect 330326 705242 330562 705478
rect 330646 705242 330882 705478
rect 330326 691718 330562 691954
rect 330646 691718 330882 691954
rect 330326 691398 330562 691634
rect 330646 691398 330882 691634
rect 330326 655718 330562 655954
rect 330646 655718 330882 655954
rect 330326 655398 330562 655634
rect 330646 655398 330882 655634
rect 330326 619718 330562 619954
rect 330646 619718 330882 619954
rect 330326 619398 330562 619634
rect 330646 619398 330882 619634
rect 330326 583718 330562 583954
rect 330646 583718 330882 583954
rect 330326 583398 330562 583634
rect 330646 583398 330882 583634
rect 330326 547718 330562 547954
rect 330646 547718 330882 547954
rect 330326 547398 330562 547634
rect 330646 547398 330882 547634
rect 330326 511718 330562 511954
rect 330646 511718 330882 511954
rect 330326 511398 330562 511634
rect 330646 511398 330882 511634
rect 330326 475718 330562 475954
rect 330646 475718 330882 475954
rect 330326 475398 330562 475634
rect 330646 475398 330882 475634
rect 330326 439718 330562 439954
rect 330646 439718 330882 439954
rect 330326 439398 330562 439634
rect 330646 439398 330882 439634
rect 330326 403718 330562 403954
rect 330646 403718 330882 403954
rect 330326 403398 330562 403634
rect 330646 403398 330882 403634
rect 330326 367718 330562 367954
rect 330646 367718 330882 367954
rect 330326 367398 330562 367634
rect 330646 367398 330882 367634
rect 330326 331718 330562 331954
rect 330646 331718 330882 331954
rect 330326 331398 330562 331634
rect 330646 331398 330882 331634
rect 330326 295718 330562 295954
rect 330646 295718 330882 295954
rect 330326 295398 330562 295634
rect 330646 295398 330882 295634
rect 330326 259718 330562 259954
rect 330646 259718 330882 259954
rect 330326 259398 330562 259634
rect 330646 259398 330882 259634
rect 330326 223718 330562 223954
rect 330646 223718 330882 223954
rect 330326 223398 330562 223634
rect 330646 223398 330882 223634
rect 330326 187718 330562 187954
rect 330646 187718 330882 187954
rect 330326 187398 330562 187634
rect 330646 187398 330882 187634
rect 334826 706522 335062 706758
rect 335146 706522 335382 706758
rect 334826 706202 335062 706438
rect 335146 706202 335382 706438
rect 334826 696218 335062 696454
rect 335146 696218 335382 696454
rect 334826 695898 335062 696134
rect 335146 695898 335382 696134
rect 334826 660218 335062 660454
rect 335146 660218 335382 660454
rect 334826 659898 335062 660134
rect 335146 659898 335382 660134
rect 334826 624218 335062 624454
rect 335146 624218 335382 624454
rect 334826 623898 335062 624134
rect 335146 623898 335382 624134
rect 334826 588218 335062 588454
rect 335146 588218 335382 588454
rect 334826 587898 335062 588134
rect 335146 587898 335382 588134
rect 334826 552218 335062 552454
rect 335146 552218 335382 552454
rect 334826 551898 335062 552134
rect 335146 551898 335382 552134
rect 334826 516218 335062 516454
rect 335146 516218 335382 516454
rect 334826 515898 335062 516134
rect 335146 515898 335382 516134
rect 334826 480218 335062 480454
rect 335146 480218 335382 480454
rect 334826 479898 335062 480134
rect 335146 479898 335382 480134
rect 334826 444218 335062 444454
rect 335146 444218 335382 444454
rect 334826 443898 335062 444134
rect 335146 443898 335382 444134
rect 334826 408218 335062 408454
rect 335146 408218 335382 408454
rect 334826 407898 335062 408134
rect 335146 407898 335382 408134
rect 334826 372218 335062 372454
rect 335146 372218 335382 372454
rect 334826 371898 335062 372134
rect 335146 371898 335382 372134
rect 334826 336218 335062 336454
rect 335146 336218 335382 336454
rect 334826 335898 335062 336134
rect 335146 335898 335382 336134
rect 334826 300218 335062 300454
rect 335146 300218 335382 300454
rect 334826 299898 335062 300134
rect 335146 299898 335382 300134
rect 334826 264218 335062 264454
rect 335146 264218 335382 264454
rect 334826 263898 335062 264134
rect 335146 263898 335382 264134
rect 334826 228218 335062 228454
rect 335146 228218 335382 228454
rect 334826 227898 335062 228134
rect 335146 227898 335382 228134
rect 334826 192218 335062 192454
rect 335146 192218 335382 192454
rect 334826 191898 335062 192134
rect 335146 191898 335382 192134
rect 339326 707482 339562 707718
rect 339646 707482 339882 707718
rect 339326 707162 339562 707398
rect 339646 707162 339882 707398
rect 339326 700718 339562 700954
rect 339646 700718 339882 700954
rect 339326 700398 339562 700634
rect 339646 700398 339882 700634
rect 339326 664718 339562 664954
rect 339646 664718 339882 664954
rect 339326 664398 339562 664634
rect 339646 664398 339882 664634
rect 339326 628718 339562 628954
rect 339646 628718 339882 628954
rect 339326 628398 339562 628634
rect 339646 628398 339882 628634
rect 339326 592718 339562 592954
rect 339646 592718 339882 592954
rect 339326 592398 339562 592634
rect 339646 592398 339882 592634
rect 339326 556718 339562 556954
rect 339646 556718 339882 556954
rect 339326 556398 339562 556634
rect 339646 556398 339882 556634
rect 339326 520718 339562 520954
rect 339646 520718 339882 520954
rect 339326 520398 339562 520634
rect 339646 520398 339882 520634
rect 339326 484718 339562 484954
rect 339646 484718 339882 484954
rect 339326 484398 339562 484634
rect 339646 484398 339882 484634
rect 339326 448718 339562 448954
rect 339646 448718 339882 448954
rect 339326 448398 339562 448634
rect 339646 448398 339882 448634
rect 339326 412718 339562 412954
rect 339646 412718 339882 412954
rect 339326 412398 339562 412634
rect 339646 412398 339882 412634
rect 343826 708442 344062 708678
rect 344146 708442 344382 708678
rect 343826 708122 344062 708358
rect 344146 708122 344382 708358
rect 343826 669218 344062 669454
rect 344146 669218 344382 669454
rect 343826 668898 344062 669134
rect 344146 668898 344382 669134
rect 343826 633218 344062 633454
rect 344146 633218 344382 633454
rect 343826 632898 344062 633134
rect 344146 632898 344382 633134
rect 343826 597218 344062 597454
rect 344146 597218 344382 597454
rect 343826 596898 344062 597134
rect 344146 596898 344382 597134
rect 343826 561218 344062 561454
rect 344146 561218 344382 561454
rect 343826 560898 344062 561134
rect 344146 560898 344382 561134
rect 343826 525218 344062 525454
rect 344146 525218 344382 525454
rect 343826 524898 344062 525134
rect 344146 524898 344382 525134
rect 343826 489218 344062 489454
rect 344146 489218 344382 489454
rect 343826 488898 344062 489134
rect 344146 488898 344382 489134
rect 343826 453218 344062 453454
rect 344146 453218 344382 453454
rect 343826 452898 344062 453134
rect 344146 452898 344382 453134
rect 343826 417218 344062 417454
rect 344146 417218 344382 417454
rect 343826 416898 344062 417134
rect 344146 416898 344382 417134
rect 339326 376718 339562 376954
rect 339646 376718 339882 376954
rect 339326 376398 339562 376634
rect 339646 376398 339882 376634
rect 339326 340718 339562 340954
rect 339646 340718 339882 340954
rect 339326 340398 339562 340634
rect 339646 340398 339882 340634
rect 339326 304718 339562 304954
rect 339646 304718 339882 304954
rect 339326 304398 339562 304634
rect 339646 304398 339882 304634
rect 339326 268718 339562 268954
rect 339646 268718 339882 268954
rect 339326 268398 339562 268634
rect 339646 268398 339882 268634
rect 339326 232718 339562 232954
rect 339646 232718 339882 232954
rect 339326 232398 339562 232634
rect 339646 232398 339882 232634
rect 339326 196718 339562 196954
rect 339646 196718 339882 196954
rect 339326 196398 339562 196634
rect 339646 196398 339882 196634
rect 339326 160718 339562 160954
rect 339646 160718 339882 160954
rect 339326 160398 339562 160634
rect 339646 160398 339882 160634
rect 279610 151718 279846 151954
rect 279610 151398 279846 151634
rect 310330 151718 310566 151954
rect 310330 151398 310566 151634
rect 341050 151718 341286 151954
rect 341050 151398 341286 151634
rect 264250 147218 264486 147454
rect 264250 146898 264486 147134
rect 294970 147218 295206 147454
rect 294970 146898 295206 147134
rect 325690 147218 325926 147454
rect 325690 146898 325926 147134
rect 279610 115718 279846 115954
rect 279610 115398 279846 115634
rect 310330 115718 310566 115954
rect 310330 115398 310566 115634
rect 341050 115718 341286 115954
rect 341050 115398 341286 115634
rect 264250 111218 264486 111454
rect 264250 110898 264486 111134
rect 294970 111218 295206 111454
rect 294970 110898 295206 111134
rect 325690 111218 325926 111454
rect 325690 110898 325926 111134
rect 348326 709402 348562 709638
rect 348646 709402 348882 709638
rect 348326 709082 348562 709318
rect 348646 709082 348882 709318
rect 348326 673718 348562 673954
rect 348646 673718 348882 673954
rect 348326 673398 348562 673634
rect 348646 673398 348882 673634
rect 348326 637718 348562 637954
rect 348646 637718 348882 637954
rect 348326 637398 348562 637634
rect 348646 637398 348882 637634
rect 348326 601718 348562 601954
rect 348646 601718 348882 601954
rect 348326 601398 348562 601634
rect 348646 601398 348882 601634
rect 348326 565718 348562 565954
rect 348646 565718 348882 565954
rect 348326 565398 348562 565634
rect 348646 565398 348882 565634
rect 348326 529718 348562 529954
rect 348646 529718 348882 529954
rect 348326 529398 348562 529634
rect 348646 529398 348882 529634
rect 348326 493718 348562 493954
rect 348646 493718 348882 493954
rect 348326 493398 348562 493634
rect 348646 493398 348882 493634
rect 348326 457718 348562 457954
rect 348646 457718 348882 457954
rect 348326 457398 348562 457634
rect 348646 457398 348882 457634
rect 348326 421718 348562 421954
rect 348646 421718 348882 421954
rect 348326 421398 348562 421634
rect 348646 421398 348882 421634
rect 348326 385718 348562 385954
rect 348646 385718 348882 385954
rect 348326 385398 348562 385634
rect 348646 385398 348882 385634
rect 343826 381218 344062 381454
rect 344146 381218 344382 381454
rect 343826 380898 344062 381134
rect 344146 380898 344382 381134
rect 343826 345218 344062 345454
rect 344146 345218 344382 345454
rect 343826 344898 344062 345134
rect 344146 344898 344382 345134
rect 343826 309218 344062 309454
rect 344146 309218 344382 309454
rect 343826 308898 344062 309134
rect 344146 308898 344382 309134
rect 343826 273218 344062 273454
rect 344146 273218 344382 273454
rect 343826 272898 344062 273134
rect 344146 272898 344382 273134
rect 343826 237218 344062 237454
rect 344146 237218 344382 237454
rect 343826 236898 344062 237134
rect 344146 236898 344382 237134
rect 343826 201218 344062 201454
rect 344146 201218 344382 201454
rect 343826 200898 344062 201134
rect 344146 200898 344382 201134
rect 343826 165218 344062 165454
rect 344146 165218 344382 165454
rect 343826 164898 344062 165134
rect 344146 164898 344382 165134
rect 262826 84218 263062 84454
rect 263146 84218 263382 84454
rect 262826 83898 263062 84134
rect 263146 83898 263382 84134
rect 262826 48218 263062 48454
rect 263146 48218 263382 48454
rect 262826 47898 263062 48134
rect 263146 47898 263382 48134
rect 262826 12218 263062 12454
rect 263146 12218 263382 12454
rect 262826 11898 263062 12134
rect 263146 11898 263382 12134
rect 258326 -1542 258562 -1306
rect 258646 -1542 258882 -1306
rect 258326 -1862 258562 -1626
rect 258646 -1862 258882 -1626
rect 262826 -2502 263062 -2266
rect 263146 -2502 263382 -2266
rect 262826 -2822 263062 -2586
rect 263146 -2822 263382 -2586
rect 267326 88718 267562 88954
rect 267646 88718 267882 88954
rect 267326 88398 267562 88634
rect 267646 88398 267882 88634
rect 267326 52718 267562 52954
rect 267646 52718 267882 52954
rect 267326 52398 267562 52634
rect 267646 52398 267882 52634
rect 267326 16718 267562 16954
rect 267646 16718 267882 16954
rect 267326 16398 267562 16634
rect 267646 16398 267882 16634
rect 267326 -3462 267562 -3226
rect 267646 -3462 267882 -3226
rect 267326 -3782 267562 -3546
rect 267646 -3782 267882 -3546
rect 271826 93218 272062 93454
rect 272146 93218 272382 93454
rect 271826 92898 272062 93134
rect 272146 92898 272382 93134
rect 271826 57218 272062 57454
rect 272146 57218 272382 57454
rect 271826 56898 272062 57134
rect 272146 56898 272382 57134
rect 271826 21218 272062 21454
rect 272146 21218 272382 21454
rect 271826 20898 272062 21134
rect 272146 20898 272382 21134
rect 271826 -4422 272062 -4186
rect 272146 -4422 272382 -4186
rect 271826 -4742 272062 -4506
rect 272146 -4742 272382 -4506
rect 276326 97718 276562 97954
rect 276646 97718 276882 97954
rect 276326 97398 276562 97634
rect 276646 97398 276882 97634
rect 276326 61718 276562 61954
rect 276646 61718 276882 61954
rect 276326 61398 276562 61634
rect 276646 61398 276882 61634
rect 276326 25718 276562 25954
rect 276646 25718 276882 25954
rect 276326 25398 276562 25634
rect 276646 25398 276882 25634
rect 276326 -5382 276562 -5146
rect 276646 -5382 276882 -5146
rect 276326 -5702 276562 -5466
rect 276646 -5702 276882 -5466
rect 280826 66218 281062 66454
rect 281146 66218 281382 66454
rect 280826 65898 281062 66134
rect 281146 65898 281382 66134
rect 280826 30218 281062 30454
rect 281146 30218 281382 30454
rect 280826 29898 281062 30134
rect 281146 29898 281382 30134
rect 280826 -6342 281062 -6106
rect 281146 -6342 281382 -6106
rect 280826 -6662 281062 -6426
rect 281146 -6662 281382 -6426
rect 285326 70718 285562 70954
rect 285646 70718 285882 70954
rect 285326 70398 285562 70634
rect 285646 70398 285882 70634
rect 285326 34718 285562 34954
rect 285646 34718 285882 34954
rect 285326 34398 285562 34634
rect 285646 34398 285882 34634
rect 285326 -7302 285562 -7066
rect 285646 -7302 285882 -7066
rect 285326 -7622 285562 -7386
rect 285646 -7622 285882 -7386
rect 289826 75218 290062 75454
rect 290146 75218 290382 75454
rect 289826 74898 290062 75134
rect 290146 74898 290382 75134
rect 289826 39218 290062 39454
rect 290146 39218 290382 39454
rect 289826 38898 290062 39134
rect 290146 38898 290382 39134
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 294326 79718 294562 79954
rect 294646 79718 294882 79954
rect 294326 79398 294562 79634
rect 294646 79398 294882 79634
rect 294326 43718 294562 43954
rect 294646 43718 294882 43954
rect 294326 43398 294562 43634
rect 294646 43398 294882 43634
rect 294326 7718 294562 7954
rect 294646 7718 294882 7954
rect 294326 7398 294562 7634
rect 294646 7398 294882 7634
rect 294326 -1542 294562 -1306
rect 294646 -1542 294882 -1306
rect 294326 -1862 294562 -1626
rect 294646 -1862 294882 -1626
rect 298826 84218 299062 84454
rect 299146 84218 299382 84454
rect 298826 83898 299062 84134
rect 299146 83898 299382 84134
rect 298826 48218 299062 48454
rect 299146 48218 299382 48454
rect 298826 47898 299062 48134
rect 299146 47898 299382 48134
rect 298826 12218 299062 12454
rect 299146 12218 299382 12454
rect 298826 11898 299062 12134
rect 299146 11898 299382 12134
rect 298826 -2502 299062 -2266
rect 299146 -2502 299382 -2266
rect 298826 -2822 299062 -2586
rect 299146 -2822 299382 -2586
rect 303326 88718 303562 88954
rect 303646 88718 303882 88954
rect 303326 88398 303562 88634
rect 303646 88398 303882 88634
rect 303326 52718 303562 52954
rect 303646 52718 303882 52954
rect 303326 52398 303562 52634
rect 303646 52398 303882 52634
rect 303326 16718 303562 16954
rect 303646 16718 303882 16954
rect 303326 16398 303562 16634
rect 303646 16398 303882 16634
rect 303326 -3462 303562 -3226
rect 303646 -3462 303882 -3226
rect 303326 -3782 303562 -3546
rect 303646 -3782 303882 -3546
rect 307826 93218 308062 93454
rect 308146 93218 308382 93454
rect 307826 92898 308062 93134
rect 308146 92898 308382 93134
rect 307826 57218 308062 57454
rect 308146 57218 308382 57454
rect 307826 56898 308062 57134
rect 308146 56898 308382 57134
rect 307826 21218 308062 21454
rect 308146 21218 308382 21454
rect 307826 20898 308062 21134
rect 308146 20898 308382 21134
rect 307826 -4422 308062 -4186
rect 308146 -4422 308382 -4186
rect 307826 -4742 308062 -4506
rect 308146 -4742 308382 -4506
rect 312326 97718 312562 97954
rect 312646 97718 312882 97954
rect 312326 97398 312562 97634
rect 312646 97398 312882 97634
rect 312326 61718 312562 61954
rect 312646 61718 312882 61954
rect 312326 61398 312562 61634
rect 312646 61398 312882 61634
rect 312326 25718 312562 25954
rect 312646 25718 312882 25954
rect 312326 25398 312562 25634
rect 312646 25398 312882 25634
rect 312326 -5382 312562 -5146
rect 312646 -5382 312882 -5146
rect 312326 -5702 312562 -5466
rect 312646 -5702 312882 -5466
rect 316826 66218 317062 66454
rect 317146 66218 317382 66454
rect 316826 65898 317062 66134
rect 317146 65898 317382 66134
rect 316826 30218 317062 30454
rect 317146 30218 317382 30454
rect 316826 29898 317062 30134
rect 317146 29898 317382 30134
rect 316826 -6342 317062 -6106
rect 317146 -6342 317382 -6106
rect 316826 -6662 317062 -6426
rect 317146 -6662 317382 -6426
rect 321326 70718 321562 70954
rect 321646 70718 321882 70954
rect 321326 70398 321562 70634
rect 321646 70398 321882 70634
rect 321326 34718 321562 34954
rect 321646 34718 321882 34954
rect 321326 34398 321562 34634
rect 321646 34398 321882 34634
rect 321326 -7302 321562 -7066
rect 321646 -7302 321882 -7066
rect 321326 -7622 321562 -7386
rect 321646 -7622 321882 -7386
rect 325826 75218 326062 75454
rect 326146 75218 326382 75454
rect 325826 74898 326062 75134
rect 326146 74898 326382 75134
rect 325826 39218 326062 39454
rect 326146 39218 326382 39454
rect 325826 38898 326062 39134
rect 326146 38898 326382 39134
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 330326 79718 330562 79954
rect 330646 79718 330882 79954
rect 330326 79398 330562 79634
rect 330646 79398 330882 79634
rect 330326 43718 330562 43954
rect 330646 43718 330882 43954
rect 330326 43398 330562 43634
rect 330646 43398 330882 43634
rect 330326 7718 330562 7954
rect 330646 7718 330882 7954
rect 330326 7398 330562 7634
rect 330646 7398 330882 7634
rect 330326 -1542 330562 -1306
rect 330646 -1542 330882 -1306
rect 330326 -1862 330562 -1626
rect 330646 -1862 330882 -1626
rect 334826 84218 335062 84454
rect 335146 84218 335382 84454
rect 334826 83898 335062 84134
rect 335146 83898 335382 84134
rect 334826 48218 335062 48454
rect 335146 48218 335382 48454
rect 334826 47898 335062 48134
rect 335146 47898 335382 48134
rect 334826 12218 335062 12454
rect 335146 12218 335382 12454
rect 334826 11898 335062 12134
rect 335146 11898 335382 12134
rect 334826 -2502 335062 -2266
rect 335146 -2502 335382 -2266
rect 334826 -2822 335062 -2586
rect 335146 -2822 335382 -2586
rect 339326 88718 339562 88954
rect 339646 88718 339882 88954
rect 339326 88398 339562 88634
rect 339646 88398 339882 88634
rect 339326 52718 339562 52954
rect 339646 52718 339882 52954
rect 339326 52398 339562 52634
rect 339646 52398 339882 52634
rect 339326 16718 339562 16954
rect 339646 16718 339882 16954
rect 339326 16398 339562 16634
rect 339646 16398 339882 16634
rect 343826 93218 344062 93454
rect 344146 93218 344382 93454
rect 343826 92898 344062 93134
rect 344146 92898 344382 93134
rect 343826 57218 344062 57454
rect 344146 57218 344382 57454
rect 343826 56898 344062 57134
rect 344146 56898 344382 57134
rect 343826 21218 344062 21454
rect 344146 21218 344382 21454
rect 343826 20898 344062 21134
rect 344146 20898 344382 21134
rect 339326 -3462 339562 -3226
rect 339646 -3462 339882 -3226
rect 339326 -3782 339562 -3546
rect 339646 -3782 339882 -3546
rect 348326 349718 348562 349954
rect 348646 349718 348882 349954
rect 348326 349398 348562 349634
rect 348646 349398 348882 349634
rect 348326 313718 348562 313954
rect 348646 313718 348882 313954
rect 348326 313398 348562 313634
rect 348646 313398 348882 313634
rect 348326 277718 348562 277954
rect 348646 277718 348882 277954
rect 348326 277398 348562 277634
rect 348646 277398 348882 277634
rect 348326 241718 348562 241954
rect 348646 241718 348882 241954
rect 348326 241398 348562 241634
rect 348646 241398 348882 241634
rect 348326 205718 348562 205954
rect 348646 205718 348882 205954
rect 348326 205398 348562 205634
rect 348646 205398 348882 205634
rect 348326 169718 348562 169954
rect 348646 169718 348882 169954
rect 348326 169398 348562 169634
rect 348646 169398 348882 169634
rect 348326 133718 348562 133954
rect 348646 133718 348882 133954
rect 348326 133398 348562 133634
rect 348646 133398 348882 133634
rect 348326 97718 348562 97954
rect 348646 97718 348882 97954
rect 348326 97398 348562 97634
rect 348646 97398 348882 97634
rect 348326 61718 348562 61954
rect 348646 61718 348882 61954
rect 348326 61398 348562 61634
rect 348646 61398 348882 61634
rect 348326 25718 348562 25954
rect 348646 25718 348882 25954
rect 348326 25398 348562 25634
rect 348646 25398 348882 25634
rect 343826 -4422 344062 -4186
rect 344146 -4422 344382 -4186
rect 343826 -4742 344062 -4506
rect 344146 -4742 344382 -4506
rect 348326 -5382 348562 -5146
rect 348646 -5382 348882 -5146
rect 348326 -5702 348562 -5466
rect 348646 -5702 348882 -5466
rect 352826 710362 353062 710598
rect 353146 710362 353382 710598
rect 352826 710042 353062 710278
rect 353146 710042 353382 710278
rect 352826 678218 353062 678454
rect 353146 678218 353382 678454
rect 352826 677898 353062 678134
rect 353146 677898 353382 678134
rect 352826 642218 353062 642454
rect 353146 642218 353382 642454
rect 352826 641898 353062 642134
rect 353146 641898 353382 642134
rect 352826 606218 353062 606454
rect 353146 606218 353382 606454
rect 352826 605898 353062 606134
rect 353146 605898 353382 606134
rect 352826 570218 353062 570454
rect 353146 570218 353382 570454
rect 352826 569898 353062 570134
rect 353146 569898 353382 570134
rect 352826 534218 353062 534454
rect 353146 534218 353382 534454
rect 352826 533898 353062 534134
rect 353146 533898 353382 534134
rect 352826 498218 353062 498454
rect 353146 498218 353382 498454
rect 352826 497898 353062 498134
rect 353146 497898 353382 498134
rect 352826 462218 353062 462454
rect 353146 462218 353382 462454
rect 352826 461898 353062 462134
rect 353146 461898 353382 462134
rect 352826 426218 353062 426454
rect 353146 426218 353382 426454
rect 352826 425898 353062 426134
rect 353146 425898 353382 426134
rect 352826 390218 353062 390454
rect 353146 390218 353382 390454
rect 352826 389898 353062 390134
rect 353146 389898 353382 390134
rect 352826 354218 353062 354454
rect 353146 354218 353382 354454
rect 352826 353898 353062 354134
rect 353146 353898 353382 354134
rect 352826 318218 353062 318454
rect 353146 318218 353382 318454
rect 352826 317898 353062 318134
rect 353146 317898 353382 318134
rect 352826 282218 353062 282454
rect 353146 282218 353382 282454
rect 352826 281898 353062 282134
rect 353146 281898 353382 282134
rect 352826 246218 353062 246454
rect 353146 246218 353382 246454
rect 352826 245898 353062 246134
rect 353146 245898 353382 246134
rect 352826 210218 353062 210454
rect 353146 210218 353382 210454
rect 352826 209898 353062 210134
rect 353146 209898 353382 210134
rect 352826 174218 353062 174454
rect 353146 174218 353382 174454
rect 352826 173898 353062 174134
rect 353146 173898 353382 174134
rect 352826 138218 353062 138454
rect 353146 138218 353382 138454
rect 352826 137898 353062 138134
rect 353146 137898 353382 138134
rect 352826 102218 353062 102454
rect 353146 102218 353382 102454
rect 352826 101898 353062 102134
rect 353146 101898 353382 102134
rect 352826 66218 353062 66454
rect 353146 66218 353382 66454
rect 352826 65898 353062 66134
rect 353146 65898 353382 66134
rect 352826 30218 353062 30454
rect 353146 30218 353382 30454
rect 352826 29898 353062 30134
rect 353146 29898 353382 30134
rect 352826 -6342 353062 -6106
rect 353146 -6342 353382 -6106
rect 352826 -6662 353062 -6426
rect 353146 -6662 353382 -6426
rect 357326 711322 357562 711558
rect 357646 711322 357882 711558
rect 357326 711002 357562 711238
rect 357646 711002 357882 711238
rect 357326 682718 357562 682954
rect 357646 682718 357882 682954
rect 357326 682398 357562 682634
rect 357646 682398 357882 682634
rect 357326 646718 357562 646954
rect 357646 646718 357882 646954
rect 357326 646398 357562 646634
rect 357646 646398 357882 646634
rect 357326 610718 357562 610954
rect 357646 610718 357882 610954
rect 357326 610398 357562 610634
rect 357646 610398 357882 610634
rect 357326 574718 357562 574954
rect 357646 574718 357882 574954
rect 357326 574398 357562 574634
rect 357646 574398 357882 574634
rect 357326 538718 357562 538954
rect 357646 538718 357882 538954
rect 357326 538398 357562 538634
rect 357646 538398 357882 538634
rect 357326 502718 357562 502954
rect 357646 502718 357882 502954
rect 357326 502398 357562 502634
rect 357646 502398 357882 502634
rect 357326 466718 357562 466954
rect 357646 466718 357882 466954
rect 357326 466398 357562 466634
rect 357646 466398 357882 466634
rect 357326 430718 357562 430954
rect 357646 430718 357882 430954
rect 357326 430398 357562 430634
rect 357646 430398 357882 430634
rect 357326 394718 357562 394954
rect 357646 394718 357882 394954
rect 357326 394398 357562 394634
rect 357646 394398 357882 394634
rect 357326 358718 357562 358954
rect 357646 358718 357882 358954
rect 357326 358398 357562 358634
rect 357646 358398 357882 358634
rect 357326 322718 357562 322954
rect 357646 322718 357882 322954
rect 357326 322398 357562 322634
rect 357646 322398 357882 322634
rect 357326 286718 357562 286954
rect 357646 286718 357882 286954
rect 357326 286398 357562 286634
rect 357646 286398 357882 286634
rect 357326 250718 357562 250954
rect 357646 250718 357882 250954
rect 357326 250398 357562 250634
rect 357646 250398 357882 250634
rect 357326 214718 357562 214954
rect 357646 214718 357882 214954
rect 357326 214398 357562 214634
rect 357646 214398 357882 214634
rect 357326 178718 357562 178954
rect 357646 178718 357882 178954
rect 357326 178398 357562 178634
rect 357646 178398 357882 178634
rect 357326 142718 357562 142954
rect 357646 142718 357882 142954
rect 357326 142398 357562 142634
rect 357646 142398 357882 142634
rect 357326 106718 357562 106954
rect 357646 106718 357882 106954
rect 357326 106398 357562 106634
rect 357646 106398 357882 106634
rect 357326 70718 357562 70954
rect 357646 70718 357882 70954
rect 357326 70398 357562 70634
rect 357646 70398 357882 70634
rect 357326 34718 357562 34954
rect 357646 34718 357882 34954
rect 357326 34398 357562 34634
rect 357646 34398 357882 34634
rect 357326 -7302 357562 -7066
rect 357646 -7302 357882 -7066
rect 357326 -7622 357562 -7386
rect 357646 -7622 357882 -7386
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 361826 651218 362062 651454
rect 362146 651218 362382 651454
rect 361826 650898 362062 651134
rect 362146 650898 362382 651134
rect 361826 615218 362062 615454
rect 362146 615218 362382 615454
rect 361826 614898 362062 615134
rect 362146 614898 362382 615134
rect 361826 579218 362062 579454
rect 362146 579218 362382 579454
rect 361826 578898 362062 579134
rect 362146 578898 362382 579134
rect 361826 543218 362062 543454
rect 362146 543218 362382 543454
rect 361826 542898 362062 543134
rect 362146 542898 362382 543134
rect 361826 507218 362062 507454
rect 362146 507218 362382 507454
rect 361826 506898 362062 507134
rect 362146 506898 362382 507134
rect 361826 471218 362062 471454
rect 362146 471218 362382 471454
rect 361826 470898 362062 471134
rect 362146 470898 362382 471134
rect 361826 435218 362062 435454
rect 362146 435218 362382 435454
rect 361826 434898 362062 435134
rect 362146 434898 362382 435134
rect 361826 399218 362062 399454
rect 362146 399218 362382 399454
rect 361826 398898 362062 399134
rect 362146 398898 362382 399134
rect 361826 363218 362062 363454
rect 362146 363218 362382 363454
rect 361826 362898 362062 363134
rect 362146 362898 362382 363134
rect 361826 327218 362062 327454
rect 362146 327218 362382 327454
rect 361826 326898 362062 327134
rect 362146 326898 362382 327134
rect 361826 291218 362062 291454
rect 362146 291218 362382 291454
rect 361826 290898 362062 291134
rect 362146 290898 362382 291134
rect 361826 255218 362062 255454
rect 362146 255218 362382 255454
rect 361826 254898 362062 255134
rect 362146 254898 362382 255134
rect 361826 219218 362062 219454
rect 362146 219218 362382 219454
rect 361826 218898 362062 219134
rect 362146 218898 362382 219134
rect 361826 183218 362062 183454
rect 362146 183218 362382 183454
rect 361826 182898 362062 183134
rect 362146 182898 362382 183134
rect 361826 147218 362062 147454
rect 362146 147218 362382 147454
rect 361826 146898 362062 147134
rect 362146 146898 362382 147134
rect 361826 111218 362062 111454
rect 362146 111218 362382 111454
rect 361826 110898 362062 111134
rect 362146 110898 362382 111134
rect 361826 75218 362062 75454
rect 362146 75218 362382 75454
rect 361826 74898 362062 75134
rect 362146 74898 362382 75134
rect 361826 39218 362062 39454
rect 362146 39218 362382 39454
rect 361826 38898 362062 39134
rect 362146 38898 362382 39134
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 366326 705562 366562 705798
rect 366646 705562 366882 705798
rect 366326 705242 366562 705478
rect 366646 705242 366882 705478
rect 366326 691718 366562 691954
rect 366646 691718 366882 691954
rect 366326 691398 366562 691634
rect 366646 691398 366882 691634
rect 366326 655718 366562 655954
rect 366646 655718 366882 655954
rect 366326 655398 366562 655634
rect 366646 655398 366882 655634
rect 366326 619718 366562 619954
rect 366646 619718 366882 619954
rect 366326 619398 366562 619634
rect 366646 619398 366882 619634
rect 366326 583718 366562 583954
rect 366646 583718 366882 583954
rect 366326 583398 366562 583634
rect 366646 583398 366882 583634
rect 366326 547718 366562 547954
rect 366646 547718 366882 547954
rect 366326 547398 366562 547634
rect 366646 547398 366882 547634
rect 366326 511718 366562 511954
rect 366646 511718 366882 511954
rect 366326 511398 366562 511634
rect 366646 511398 366882 511634
rect 366326 475718 366562 475954
rect 366646 475718 366882 475954
rect 366326 475398 366562 475634
rect 366646 475398 366882 475634
rect 366326 439718 366562 439954
rect 366646 439718 366882 439954
rect 366326 439398 366562 439634
rect 366646 439398 366882 439634
rect 366326 403718 366562 403954
rect 366646 403718 366882 403954
rect 366326 403398 366562 403634
rect 366646 403398 366882 403634
rect 366326 367718 366562 367954
rect 366646 367718 366882 367954
rect 366326 367398 366562 367634
rect 366646 367398 366882 367634
rect 366326 331718 366562 331954
rect 366646 331718 366882 331954
rect 366326 331398 366562 331634
rect 366646 331398 366882 331634
rect 366326 295718 366562 295954
rect 366646 295718 366882 295954
rect 366326 295398 366562 295634
rect 366646 295398 366882 295634
rect 366326 259718 366562 259954
rect 366646 259718 366882 259954
rect 366326 259398 366562 259634
rect 366646 259398 366882 259634
rect 366326 223718 366562 223954
rect 366646 223718 366882 223954
rect 366326 223398 366562 223634
rect 366646 223398 366882 223634
rect 366326 187718 366562 187954
rect 366646 187718 366882 187954
rect 366326 187398 366562 187634
rect 366646 187398 366882 187634
rect 366326 151718 366562 151954
rect 366646 151718 366882 151954
rect 366326 151398 366562 151634
rect 366646 151398 366882 151634
rect 366326 115718 366562 115954
rect 366646 115718 366882 115954
rect 366326 115398 366562 115634
rect 366646 115398 366882 115634
rect 366326 79718 366562 79954
rect 366646 79718 366882 79954
rect 366326 79398 366562 79634
rect 366646 79398 366882 79634
rect 366326 43718 366562 43954
rect 366646 43718 366882 43954
rect 366326 43398 366562 43634
rect 366646 43398 366882 43634
rect 366326 7718 366562 7954
rect 366646 7718 366882 7954
rect 366326 7398 366562 7634
rect 366646 7398 366882 7634
rect 366326 -1542 366562 -1306
rect 366646 -1542 366882 -1306
rect 366326 -1862 366562 -1626
rect 366646 -1862 366882 -1626
rect 370826 706522 371062 706758
rect 371146 706522 371382 706758
rect 370826 706202 371062 706438
rect 371146 706202 371382 706438
rect 370826 696218 371062 696454
rect 371146 696218 371382 696454
rect 370826 695898 371062 696134
rect 371146 695898 371382 696134
rect 370826 660218 371062 660454
rect 371146 660218 371382 660454
rect 370826 659898 371062 660134
rect 371146 659898 371382 660134
rect 370826 624218 371062 624454
rect 371146 624218 371382 624454
rect 370826 623898 371062 624134
rect 371146 623898 371382 624134
rect 370826 588218 371062 588454
rect 371146 588218 371382 588454
rect 370826 587898 371062 588134
rect 371146 587898 371382 588134
rect 370826 552218 371062 552454
rect 371146 552218 371382 552454
rect 370826 551898 371062 552134
rect 371146 551898 371382 552134
rect 370826 516218 371062 516454
rect 371146 516218 371382 516454
rect 370826 515898 371062 516134
rect 371146 515898 371382 516134
rect 370826 480218 371062 480454
rect 371146 480218 371382 480454
rect 370826 479898 371062 480134
rect 371146 479898 371382 480134
rect 370826 444218 371062 444454
rect 371146 444218 371382 444454
rect 370826 443898 371062 444134
rect 371146 443898 371382 444134
rect 370826 408218 371062 408454
rect 371146 408218 371382 408454
rect 370826 407898 371062 408134
rect 371146 407898 371382 408134
rect 370826 372218 371062 372454
rect 371146 372218 371382 372454
rect 370826 371898 371062 372134
rect 371146 371898 371382 372134
rect 370826 336218 371062 336454
rect 371146 336218 371382 336454
rect 370826 335898 371062 336134
rect 371146 335898 371382 336134
rect 370826 300218 371062 300454
rect 371146 300218 371382 300454
rect 370826 299898 371062 300134
rect 371146 299898 371382 300134
rect 370826 264218 371062 264454
rect 371146 264218 371382 264454
rect 370826 263898 371062 264134
rect 371146 263898 371382 264134
rect 370826 228218 371062 228454
rect 371146 228218 371382 228454
rect 370826 227898 371062 228134
rect 371146 227898 371382 228134
rect 370826 192218 371062 192454
rect 371146 192218 371382 192454
rect 370826 191898 371062 192134
rect 371146 191898 371382 192134
rect 370826 156218 371062 156454
rect 371146 156218 371382 156454
rect 370826 155898 371062 156134
rect 371146 155898 371382 156134
rect 370826 120218 371062 120454
rect 371146 120218 371382 120454
rect 370826 119898 371062 120134
rect 371146 119898 371382 120134
rect 370826 84218 371062 84454
rect 371146 84218 371382 84454
rect 370826 83898 371062 84134
rect 371146 83898 371382 84134
rect 370826 48218 371062 48454
rect 371146 48218 371382 48454
rect 370826 47898 371062 48134
rect 371146 47898 371382 48134
rect 370826 12218 371062 12454
rect 371146 12218 371382 12454
rect 370826 11898 371062 12134
rect 371146 11898 371382 12134
rect 370826 -2502 371062 -2266
rect 371146 -2502 371382 -2266
rect 370826 -2822 371062 -2586
rect 371146 -2822 371382 -2586
rect 375326 707482 375562 707718
rect 375646 707482 375882 707718
rect 375326 707162 375562 707398
rect 375646 707162 375882 707398
rect 375326 700718 375562 700954
rect 375646 700718 375882 700954
rect 375326 700398 375562 700634
rect 375646 700398 375882 700634
rect 375326 664718 375562 664954
rect 375646 664718 375882 664954
rect 375326 664398 375562 664634
rect 375646 664398 375882 664634
rect 375326 628718 375562 628954
rect 375646 628718 375882 628954
rect 375326 628398 375562 628634
rect 375646 628398 375882 628634
rect 375326 592718 375562 592954
rect 375646 592718 375882 592954
rect 375326 592398 375562 592634
rect 375646 592398 375882 592634
rect 379826 708442 380062 708678
rect 380146 708442 380382 708678
rect 379826 708122 380062 708358
rect 380146 708122 380382 708358
rect 379826 669218 380062 669454
rect 380146 669218 380382 669454
rect 379826 668898 380062 669134
rect 380146 668898 380382 669134
rect 379826 633218 380062 633454
rect 380146 633218 380382 633454
rect 379826 632898 380062 633134
rect 380146 632898 380382 633134
rect 379826 597218 380062 597454
rect 380146 597218 380382 597454
rect 379826 596898 380062 597134
rect 380146 596898 380382 597134
rect 384326 709402 384562 709638
rect 384646 709402 384882 709638
rect 384326 709082 384562 709318
rect 384646 709082 384882 709318
rect 384326 673718 384562 673954
rect 384646 673718 384882 673954
rect 384326 673398 384562 673634
rect 384646 673398 384882 673634
rect 384326 637718 384562 637954
rect 384646 637718 384882 637954
rect 384326 637398 384562 637634
rect 384646 637398 384882 637634
rect 384326 601718 384562 601954
rect 384646 601718 384882 601954
rect 384326 601398 384562 601634
rect 384646 601398 384882 601634
rect 388826 710362 389062 710598
rect 389146 710362 389382 710598
rect 388826 710042 389062 710278
rect 389146 710042 389382 710278
rect 388826 678218 389062 678454
rect 389146 678218 389382 678454
rect 388826 677898 389062 678134
rect 389146 677898 389382 678134
rect 388826 642218 389062 642454
rect 389146 642218 389382 642454
rect 388826 641898 389062 642134
rect 389146 641898 389382 642134
rect 388826 606218 389062 606454
rect 389146 606218 389382 606454
rect 388826 605898 389062 606134
rect 389146 605898 389382 606134
rect 393326 711322 393562 711558
rect 393646 711322 393882 711558
rect 393326 711002 393562 711238
rect 393646 711002 393882 711238
rect 393326 682718 393562 682954
rect 393646 682718 393882 682954
rect 393326 682398 393562 682634
rect 393646 682398 393882 682634
rect 393326 646718 393562 646954
rect 393646 646718 393882 646954
rect 393326 646398 393562 646634
rect 393646 646398 393882 646634
rect 393326 610718 393562 610954
rect 393646 610718 393882 610954
rect 393326 610398 393562 610634
rect 393646 610398 393882 610634
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 397826 651218 398062 651454
rect 398146 651218 398382 651454
rect 397826 650898 398062 651134
rect 398146 650898 398382 651134
rect 397826 615218 398062 615454
rect 398146 615218 398382 615454
rect 397826 614898 398062 615134
rect 398146 614898 398382 615134
rect 402326 705562 402562 705798
rect 402646 705562 402882 705798
rect 402326 705242 402562 705478
rect 402646 705242 402882 705478
rect 402326 691718 402562 691954
rect 402646 691718 402882 691954
rect 402326 691398 402562 691634
rect 402646 691398 402882 691634
rect 402326 655718 402562 655954
rect 402646 655718 402882 655954
rect 402326 655398 402562 655634
rect 402646 655398 402882 655634
rect 402326 619718 402562 619954
rect 402646 619718 402882 619954
rect 402326 619398 402562 619634
rect 402646 619398 402882 619634
rect 406826 706522 407062 706758
rect 407146 706522 407382 706758
rect 406826 706202 407062 706438
rect 407146 706202 407382 706438
rect 406826 696218 407062 696454
rect 407146 696218 407382 696454
rect 406826 695898 407062 696134
rect 407146 695898 407382 696134
rect 406826 660218 407062 660454
rect 407146 660218 407382 660454
rect 406826 659898 407062 660134
rect 407146 659898 407382 660134
rect 406826 624218 407062 624454
rect 407146 624218 407382 624454
rect 406826 623898 407062 624134
rect 407146 623898 407382 624134
rect 411326 707482 411562 707718
rect 411646 707482 411882 707718
rect 411326 707162 411562 707398
rect 411646 707162 411882 707398
rect 411326 700718 411562 700954
rect 411646 700718 411882 700954
rect 411326 700398 411562 700634
rect 411646 700398 411882 700634
rect 411326 664718 411562 664954
rect 411646 664718 411882 664954
rect 411326 664398 411562 664634
rect 411646 664398 411882 664634
rect 411326 628718 411562 628954
rect 411646 628718 411882 628954
rect 411326 628398 411562 628634
rect 411646 628398 411882 628634
rect 411326 592718 411562 592954
rect 411646 592718 411882 592954
rect 411326 592398 411562 592634
rect 411646 592398 411882 592634
rect 415826 708442 416062 708678
rect 416146 708442 416382 708678
rect 415826 708122 416062 708358
rect 416146 708122 416382 708358
rect 415826 669218 416062 669454
rect 416146 669218 416382 669454
rect 415826 668898 416062 669134
rect 416146 668898 416382 669134
rect 415826 633218 416062 633454
rect 416146 633218 416382 633454
rect 415826 632898 416062 633134
rect 416146 632898 416382 633134
rect 415826 597218 416062 597454
rect 416146 597218 416382 597454
rect 415826 596898 416062 597134
rect 416146 596898 416382 597134
rect 420326 709402 420562 709638
rect 420646 709402 420882 709638
rect 420326 709082 420562 709318
rect 420646 709082 420882 709318
rect 420326 673718 420562 673954
rect 420646 673718 420882 673954
rect 420326 673398 420562 673634
rect 420646 673398 420882 673634
rect 420326 637718 420562 637954
rect 420646 637718 420882 637954
rect 420326 637398 420562 637634
rect 420646 637398 420882 637634
rect 420326 601718 420562 601954
rect 420646 601718 420882 601954
rect 420326 601398 420562 601634
rect 420646 601398 420882 601634
rect 424826 710362 425062 710598
rect 425146 710362 425382 710598
rect 424826 710042 425062 710278
rect 425146 710042 425382 710278
rect 424826 678218 425062 678454
rect 425146 678218 425382 678454
rect 424826 677898 425062 678134
rect 425146 677898 425382 678134
rect 424826 642218 425062 642454
rect 425146 642218 425382 642454
rect 424826 641898 425062 642134
rect 425146 641898 425382 642134
rect 424826 606218 425062 606454
rect 425146 606218 425382 606454
rect 424826 605898 425062 606134
rect 425146 605898 425382 606134
rect 429326 711322 429562 711558
rect 429646 711322 429882 711558
rect 429326 711002 429562 711238
rect 429646 711002 429882 711238
rect 429326 682718 429562 682954
rect 429646 682718 429882 682954
rect 429326 682398 429562 682634
rect 429646 682398 429882 682634
rect 429326 646718 429562 646954
rect 429646 646718 429882 646954
rect 429326 646398 429562 646634
rect 429646 646398 429882 646634
rect 429326 610718 429562 610954
rect 429646 610718 429882 610954
rect 429326 610398 429562 610634
rect 429646 610398 429882 610634
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 433826 651218 434062 651454
rect 434146 651218 434382 651454
rect 433826 650898 434062 651134
rect 434146 650898 434382 651134
rect 433826 615218 434062 615454
rect 434146 615218 434382 615454
rect 433826 614898 434062 615134
rect 434146 614898 434382 615134
rect 438326 705562 438562 705798
rect 438646 705562 438882 705798
rect 438326 705242 438562 705478
rect 438646 705242 438882 705478
rect 438326 691718 438562 691954
rect 438646 691718 438882 691954
rect 438326 691398 438562 691634
rect 438646 691398 438882 691634
rect 438326 655718 438562 655954
rect 438646 655718 438882 655954
rect 438326 655398 438562 655634
rect 438646 655398 438882 655634
rect 438326 619718 438562 619954
rect 438646 619718 438882 619954
rect 438326 619398 438562 619634
rect 438646 619398 438882 619634
rect 442826 706522 443062 706758
rect 443146 706522 443382 706758
rect 442826 706202 443062 706438
rect 443146 706202 443382 706438
rect 442826 696218 443062 696454
rect 443146 696218 443382 696454
rect 442826 695898 443062 696134
rect 443146 695898 443382 696134
rect 442826 660218 443062 660454
rect 443146 660218 443382 660454
rect 442826 659898 443062 660134
rect 443146 659898 443382 660134
rect 442826 624218 443062 624454
rect 443146 624218 443382 624454
rect 442826 623898 443062 624134
rect 443146 623898 443382 624134
rect 447326 707482 447562 707718
rect 447646 707482 447882 707718
rect 447326 707162 447562 707398
rect 447646 707162 447882 707398
rect 447326 700718 447562 700954
rect 447646 700718 447882 700954
rect 447326 700398 447562 700634
rect 447646 700398 447882 700634
rect 447326 664718 447562 664954
rect 447646 664718 447882 664954
rect 447326 664398 447562 664634
rect 447646 664398 447882 664634
rect 447326 628718 447562 628954
rect 447646 628718 447882 628954
rect 447326 628398 447562 628634
rect 447646 628398 447882 628634
rect 447326 592718 447562 592954
rect 447646 592718 447882 592954
rect 447326 592398 447562 592634
rect 447646 592398 447882 592634
rect 451826 708442 452062 708678
rect 452146 708442 452382 708678
rect 451826 708122 452062 708358
rect 452146 708122 452382 708358
rect 451826 669218 452062 669454
rect 452146 669218 452382 669454
rect 451826 668898 452062 669134
rect 452146 668898 452382 669134
rect 451826 633218 452062 633454
rect 452146 633218 452382 633454
rect 451826 632898 452062 633134
rect 452146 632898 452382 633134
rect 451826 597218 452062 597454
rect 452146 597218 452382 597454
rect 451826 596898 452062 597134
rect 452146 596898 452382 597134
rect 456326 709402 456562 709638
rect 456646 709402 456882 709638
rect 456326 709082 456562 709318
rect 456646 709082 456882 709318
rect 456326 673718 456562 673954
rect 456646 673718 456882 673954
rect 456326 673398 456562 673634
rect 456646 673398 456882 673634
rect 456326 637718 456562 637954
rect 456646 637718 456882 637954
rect 456326 637398 456562 637634
rect 456646 637398 456882 637634
rect 456326 601718 456562 601954
rect 456646 601718 456882 601954
rect 456326 601398 456562 601634
rect 456646 601398 456882 601634
rect 460826 710362 461062 710598
rect 461146 710362 461382 710598
rect 460826 710042 461062 710278
rect 461146 710042 461382 710278
rect 460826 678218 461062 678454
rect 461146 678218 461382 678454
rect 460826 677898 461062 678134
rect 461146 677898 461382 678134
rect 460826 642218 461062 642454
rect 461146 642218 461382 642454
rect 460826 641898 461062 642134
rect 461146 641898 461382 642134
rect 460826 606218 461062 606454
rect 461146 606218 461382 606454
rect 460826 605898 461062 606134
rect 461146 605898 461382 606134
rect 465326 711322 465562 711558
rect 465646 711322 465882 711558
rect 465326 711002 465562 711238
rect 465646 711002 465882 711238
rect 465326 682718 465562 682954
rect 465646 682718 465882 682954
rect 465326 682398 465562 682634
rect 465646 682398 465882 682634
rect 465326 646718 465562 646954
rect 465646 646718 465882 646954
rect 465326 646398 465562 646634
rect 465646 646398 465882 646634
rect 465326 610718 465562 610954
rect 465646 610718 465882 610954
rect 465326 610398 465562 610634
rect 465646 610398 465882 610634
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 469826 651218 470062 651454
rect 470146 651218 470382 651454
rect 469826 650898 470062 651134
rect 470146 650898 470382 651134
rect 469826 615218 470062 615454
rect 470146 615218 470382 615454
rect 469826 614898 470062 615134
rect 470146 614898 470382 615134
rect 474326 705562 474562 705798
rect 474646 705562 474882 705798
rect 474326 705242 474562 705478
rect 474646 705242 474882 705478
rect 474326 691718 474562 691954
rect 474646 691718 474882 691954
rect 474326 691398 474562 691634
rect 474646 691398 474882 691634
rect 474326 655718 474562 655954
rect 474646 655718 474882 655954
rect 474326 655398 474562 655634
rect 474646 655398 474882 655634
rect 474326 619718 474562 619954
rect 474646 619718 474882 619954
rect 474326 619398 474562 619634
rect 474646 619398 474882 619634
rect 380328 583718 380564 583954
rect 380328 583398 380564 583634
rect 470496 583718 470732 583954
rect 470496 583398 470732 583634
rect 474326 583718 474562 583954
rect 474646 583718 474882 583954
rect 474326 583398 474562 583634
rect 474646 583398 474882 583634
rect 381008 579218 381244 579454
rect 381008 578898 381244 579134
rect 469816 579218 470052 579454
rect 469816 578898 470052 579134
rect 375326 556718 375562 556954
rect 375646 556718 375882 556954
rect 375326 556398 375562 556634
rect 375646 556398 375882 556634
rect 380328 547718 380564 547954
rect 380328 547398 380564 547634
rect 470496 547718 470732 547954
rect 470496 547398 470732 547634
rect 474326 547718 474562 547954
rect 474646 547718 474882 547954
rect 474326 547398 474562 547634
rect 474646 547398 474882 547634
rect 381008 543218 381244 543454
rect 381008 542898 381244 543134
rect 469816 543218 470052 543454
rect 469816 542898 470052 543134
rect 375326 520718 375562 520954
rect 375646 520718 375882 520954
rect 375326 520398 375562 520634
rect 375646 520398 375882 520634
rect 380328 511718 380564 511954
rect 380328 511398 380564 511634
rect 470496 511718 470732 511954
rect 470496 511398 470732 511634
rect 474326 511718 474562 511954
rect 474646 511718 474882 511954
rect 474326 511398 474562 511634
rect 474646 511398 474882 511634
rect 381008 507218 381244 507454
rect 381008 506898 381244 507134
rect 469816 507218 470052 507454
rect 469816 506898 470052 507134
rect 375326 484718 375562 484954
rect 375646 484718 375882 484954
rect 375326 484398 375562 484634
rect 375646 484398 375882 484634
rect 375326 448718 375562 448954
rect 375646 448718 375882 448954
rect 375326 448398 375562 448634
rect 375646 448398 375882 448634
rect 375326 412718 375562 412954
rect 375646 412718 375882 412954
rect 375326 412398 375562 412634
rect 375646 412398 375882 412634
rect 375326 376718 375562 376954
rect 375646 376718 375882 376954
rect 375326 376398 375562 376634
rect 375646 376398 375882 376634
rect 375326 340718 375562 340954
rect 375646 340718 375882 340954
rect 375326 340398 375562 340634
rect 375646 340398 375882 340634
rect 375326 304718 375562 304954
rect 375646 304718 375882 304954
rect 375326 304398 375562 304634
rect 375646 304398 375882 304634
rect 375326 268718 375562 268954
rect 375646 268718 375882 268954
rect 375326 268398 375562 268634
rect 375646 268398 375882 268634
rect 375326 232718 375562 232954
rect 375646 232718 375882 232954
rect 375326 232398 375562 232634
rect 375646 232398 375882 232634
rect 375326 196718 375562 196954
rect 375646 196718 375882 196954
rect 375326 196398 375562 196634
rect 375646 196398 375882 196634
rect 375326 160718 375562 160954
rect 375646 160718 375882 160954
rect 375326 160398 375562 160634
rect 375646 160398 375882 160634
rect 375326 124718 375562 124954
rect 375646 124718 375882 124954
rect 375326 124398 375562 124634
rect 375646 124398 375882 124634
rect 375326 88718 375562 88954
rect 375646 88718 375882 88954
rect 375326 88398 375562 88634
rect 375646 88398 375882 88634
rect 375326 52718 375562 52954
rect 375646 52718 375882 52954
rect 375326 52398 375562 52634
rect 375646 52398 375882 52634
rect 375326 16718 375562 16954
rect 375646 16718 375882 16954
rect 375326 16398 375562 16634
rect 375646 16398 375882 16634
rect 375326 -3462 375562 -3226
rect 375646 -3462 375882 -3226
rect 375326 -3782 375562 -3546
rect 375646 -3782 375882 -3546
rect 379826 489218 380062 489454
rect 380146 489218 380382 489454
rect 379826 488898 380062 489134
rect 380146 488898 380382 489134
rect 379826 453218 380062 453454
rect 380146 453218 380382 453454
rect 379826 452898 380062 453134
rect 380146 452898 380382 453134
rect 379826 417218 380062 417454
rect 380146 417218 380382 417454
rect 379826 416898 380062 417134
rect 380146 416898 380382 417134
rect 379826 381218 380062 381454
rect 380146 381218 380382 381454
rect 379826 380898 380062 381134
rect 380146 380898 380382 381134
rect 379826 345218 380062 345454
rect 380146 345218 380382 345454
rect 379826 344898 380062 345134
rect 380146 344898 380382 345134
rect 379826 309218 380062 309454
rect 380146 309218 380382 309454
rect 379826 308898 380062 309134
rect 380146 308898 380382 309134
rect 379826 273218 380062 273454
rect 380146 273218 380382 273454
rect 379826 272898 380062 273134
rect 380146 272898 380382 273134
rect 379826 237218 380062 237454
rect 380146 237218 380382 237454
rect 379826 236898 380062 237134
rect 380146 236898 380382 237134
rect 379826 201218 380062 201454
rect 380146 201218 380382 201454
rect 379826 200898 380062 201134
rect 380146 200898 380382 201134
rect 379826 165218 380062 165454
rect 380146 165218 380382 165454
rect 379826 164898 380062 165134
rect 380146 164898 380382 165134
rect 379826 129218 380062 129454
rect 380146 129218 380382 129454
rect 379826 128898 380062 129134
rect 380146 128898 380382 129134
rect 379826 93218 380062 93454
rect 380146 93218 380382 93454
rect 379826 92898 380062 93134
rect 380146 92898 380382 93134
rect 379826 57218 380062 57454
rect 380146 57218 380382 57454
rect 379826 56898 380062 57134
rect 380146 56898 380382 57134
rect 379826 21218 380062 21454
rect 380146 21218 380382 21454
rect 379826 20898 380062 21134
rect 380146 20898 380382 21134
rect 379826 -4422 380062 -4186
rect 380146 -4422 380382 -4186
rect 379826 -4742 380062 -4506
rect 380146 -4742 380382 -4506
rect 384326 493718 384562 493954
rect 384646 493718 384882 493954
rect 384326 493398 384562 493634
rect 384646 493398 384882 493634
rect 384326 457718 384562 457954
rect 384646 457718 384882 457954
rect 384326 457398 384562 457634
rect 384646 457398 384882 457634
rect 384326 421718 384562 421954
rect 384646 421718 384882 421954
rect 384326 421398 384562 421634
rect 384646 421398 384882 421634
rect 384326 385718 384562 385954
rect 384646 385718 384882 385954
rect 384326 385398 384562 385634
rect 384646 385398 384882 385634
rect 384326 349718 384562 349954
rect 384646 349718 384882 349954
rect 384326 349398 384562 349634
rect 384646 349398 384882 349634
rect 384326 313718 384562 313954
rect 384646 313718 384882 313954
rect 384326 313398 384562 313634
rect 384646 313398 384882 313634
rect 384326 277718 384562 277954
rect 384646 277718 384882 277954
rect 384326 277398 384562 277634
rect 384646 277398 384882 277634
rect 384326 241718 384562 241954
rect 384646 241718 384882 241954
rect 384326 241398 384562 241634
rect 384646 241398 384882 241634
rect 384326 205718 384562 205954
rect 384646 205718 384882 205954
rect 384326 205398 384562 205634
rect 384646 205398 384882 205634
rect 384326 169718 384562 169954
rect 384646 169718 384882 169954
rect 384326 169398 384562 169634
rect 384646 169398 384882 169634
rect 384326 133718 384562 133954
rect 384646 133718 384882 133954
rect 384326 133398 384562 133634
rect 384646 133398 384882 133634
rect 384326 97718 384562 97954
rect 384646 97718 384882 97954
rect 384326 97398 384562 97634
rect 384646 97398 384882 97634
rect 384326 61718 384562 61954
rect 384646 61718 384882 61954
rect 384326 61398 384562 61634
rect 384646 61398 384882 61634
rect 384326 25718 384562 25954
rect 384646 25718 384882 25954
rect 384326 25398 384562 25634
rect 384646 25398 384882 25634
rect 384326 -5382 384562 -5146
rect 384646 -5382 384882 -5146
rect 384326 -5702 384562 -5466
rect 384646 -5702 384882 -5466
rect 388826 462218 389062 462454
rect 389146 462218 389382 462454
rect 388826 461898 389062 462134
rect 389146 461898 389382 462134
rect 388826 426218 389062 426454
rect 389146 426218 389382 426454
rect 388826 425898 389062 426134
rect 389146 425898 389382 426134
rect 388826 390218 389062 390454
rect 389146 390218 389382 390454
rect 388826 389898 389062 390134
rect 389146 389898 389382 390134
rect 388826 354218 389062 354454
rect 389146 354218 389382 354454
rect 388826 353898 389062 354134
rect 389146 353898 389382 354134
rect 388826 318218 389062 318454
rect 389146 318218 389382 318454
rect 388826 317898 389062 318134
rect 389146 317898 389382 318134
rect 388826 282218 389062 282454
rect 389146 282218 389382 282454
rect 388826 281898 389062 282134
rect 389146 281898 389382 282134
rect 388826 246218 389062 246454
rect 389146 246218 389382 246454
rect 388826 245898 389062 246134
rect 389146 245898 389382 246134
rect 388826 210218 389062 210454
rect 389146 210218 389382 210454
rect 388826 209898 389062 210134
rect 389146 209898 389382 210134
rect 388826 174218 389062 174454
rect 389146 174218 389382 174454
rect 388826 173898 389062 174134
rect 389146 173898 389382 174134
rect 388826 138218 389062 138454
rect 389146 138218 389382 138454
rect 388826 137898 389062 138134
rect 389146 137898 389382 138134
rect 388826 102218 389062 102454
rect 389146 102218 389382 102454
rect 388826 101898 389062 102134
rect 389146 101898 389382 102134
rect 388826 66218 389062 66454
rect 389146 66218 389382 66454
rect 388826 65898 389062 66134
rect 389146 65898 389382 66134
rect 388826 30218 389062 30454
rect 389146 30218 389382 30454
rect 388826 29898 389062 30134
rect 389146 29898 389382 30134
rect 388826 -6342 389062 -6106
rect 389146 -6342 389382 -6106
rect 388826 -6662 389062 -6426
rect 389146 -6662 389382 -6426
rect 393326 466718 393562 466954
rect 393646 466718 393882 466954
rect 393326 466398 393562 466634
rect 393646 466398 393882 466634
rect 393326 430718 393562 430954
rect 393646 430718 393882 430954
rect 393326 430398 393562 430634
rect 393646 430398 393882 430634
rect 393326 394718 393562 394954
rect 393646 394718 393882 394954
rect 393326 394398 393562 394634
rect 393646 394398 393882 394634
rect 393326 358718 393562 358954
rect 393646 358718 393882 358954
rect 393326 358398 393562 358634
rect 393646 358398 393882 358634
rect 393326 322718 393562 322954
rect 393646 322718 393882 322954
rect 393326 322398 393562 322634
rect 393646 322398 393882 322634
rect 393326 286718 393562 286954
rect 393646 286718 393882 286954
rect 393326 286398 393562 286634
rect 393646 286398 393882 286634
rect 393326 250718 393562 250954
rect 393646 250718 393882 250954
rect 393326 250398 393562 250634
rect 393646 250398 393882 250634
rect 393326 214718 393562 214954
rect 393646 214718 393882 214954
rect 393326 214398 393562 214634
rect 393646 214398 393882 214634
rect 393326 178718 393562 178954
rect 393646 178718 393882 178954
rect 393326 178398 393562 178634
rect 393646 178398 393882 178634
rect 393326 142718 393562 142954
rect 393646 142718 393882 142954
rect 393326 142398 393562 142634
rect 393646 142398 393882 142634
rect 393326 106718 393562 106954
rect 393646 106718 393882 106954
rect 393326 106398 393562 106634
rect 393646 106398 393882 106634
rect 393326 70718 393562 70954
rect 393646 70718 393882 70954
rect 393326 70398 393562 70634
rect 393646 70398 393882 70634
rect 393326 34718 393562 34954
rect 393646 34718 393882 34954
rect 393326 34398 393562 34634
rect 393646 34398 393882 34634
rect 393326 -7302 393562 -7066
rect 393646 -7302 393882 -7066
rect 393326 -7622 393562 -7386
rect 393646 -7622 393882 -7386
rect 397826 471218 398062 471454
rect 398146 471218 398382 471454
rect 397826 470898 398062 471134
rect 398146 470898 398382 471134
rect 397826 435218 398062 435454
rect 398146 435218 398382 435454
rect 397826 434898 398062 435134
rect 398146 434898 398382 435134
rect 397826 399218 398062 399454
rect 398146 399218 398382 399454
rect 397826 398898 398062 399134
rect 398146 398898 398382 399134
rect 397826 363218 398062 363454
rect 398146 363218 398382 363454
rect 397826 362898 398062 363134
rect 398146 362898 398382 363134
rect 397826 327218 398062 327454
rect 398146 327218 398382 327454
rect 397826 326898 398062 327134
rect 398146 326898 398382 327134
rect 397826 291218 398062 291454
rect 398146 291218 398382 291454
rect 397826 290898 398062 291134
rect 398146 290898 398382 291134
rect 397826 255218 398062 255454
rect 398146 255218 398382 255454
rect 397826 254898 398062 255134
rect 398146 254898 398382 255134
rect 397826 219218 398062 219454
rect 398146 219218 398382 219454
rect 397826 218898 398062 219134
rect 398146 218898 398382 219134
rect 397826 183218 398062 183454
rect 398146 183218 398382 183454
rect 397826 182898 398062 183134
rect 398146 182898 398382 183134
rect 397826 147218 398062 147454
rect 398146 147218 398382 147454
rect 397826 146898 398062 147134
rect 398146 146898 398382 147134
rect 397826 111218 398062 111454
rect 398146 111218 398382 111454
rect 397826 110898 398062 111134
rect 398146 110898 398382 111134
rect 397826 75218 398062 75454
rect 398146 75218 398382 75454
rect 397826 74898 398062 75134
rect 398146 74898 398382 75134
rect 397826 39218 398062 39454
rect 398146 39218 398382 39454
rect 397826 38898 398062 39134
rect 398146 38898 398382 39134
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 402326 475718 402562 475954
rect 402646 475718 402882 475954
rect 402326 475398 402562 475634
rect 402646 475398 402882 475634
rect 402326 439718 402562 439954
rect 402646 439718 402882 439954
rect 402326 439398 402562 439634
rect 402646 439398 402882 439634
rect 402326 403718 402562 403954
rect 402646 403718 402882 403954
rect 402326 403398 402562 403634
rect 402646 403398 402882 403634
rect 402326 367718 402562 367954
rect 402646 367718 402882 367954
rect 402326 367398 402562 367634
rect 402646 367398 402882 367634
rect 402326 331718 402562 331954
rect 402646 331718 402882 331954
rect 402326 331398 402562 331634
rect 402646 331398 402882 331634
rect 402326 295718 402562 295954
rect 402646 295718 402882 295954
rect 402326 295398 402562 295634
rect 402646 295398 402882 295634
rect 402326 259718 402562 259954
rect 402646 259718 402882 259954
rect 402326 259398 402562 259634
rect 402646 259398 402882 259634
rect 402326 223718 402562 223954
rect 402646 223718 402882 223954
rect 402326 223398 402562 223634
rect 402646 223398 402882 223634
rect 402326 187718 402562 187954
rect 402646 187718 402882 187954
rect 402326 187398 402562 187634
rect 402646 187398 402882 187634
rect 402326 151718 402562 151954
rect 402646 151718 402882 151954
rect 402326 151398 402562 151634
rect 402646 151398 402882 151634
rect 402326 115718 402562 115954
rect 402646 115718 402882 115954
rect 402326 115398 402562 115634
rect 402646 115398 402882 115634
rect 402326 79718 402562 79954
rect 402646 79718 402882 79954
rect 402326 79398 402562 79634
rect 402646 79398 402882 79634
rect 402326 43718 402562 43954
rect 402646 43718 402882 43954
rect 402326 43398 402562 43634
rect 402646 43398 402882 43634
rect 402326 7718 402562 7954
rect 402646 7718 402882 7954
rect 402326 7398 402562 7634
rect 402646 7398 402882 7634
rect 402326 -1542 402562 -1306
rect 402646 -1542 402882 -1306
rect 402326 -1862 402562 -1626
rect 402646 -1862 402882 -1626
rect 406826 480218 407062 480454
rect 407146 480218 407382 480454
rect 406826 479898 407062 480134
rect 407146 479898 407382 480134
rect 406826 444218 407062 444454
rect 407146 444218 407382 444454
rect 406826 443898 407062 444134
rect 407146 443898 407382 444134
rect 406826 408218 407062 408454
rect 407146 408218 407382 408454
rect 406826 407898 407062 408134
rect 407146 407898 407382 408134
rect 406826 372218 407062 372454
rect 407146 372218 407382 372454
rect 406826 371898 407062 372134
rect 407146 371898 407382 372134
rect 406826 336218 407062 336454
rect 407146 336218 407382 336454
rect 406826 335898 407062 336134
rect 407146 335898 407382 336134
rect 406826 300218 407062 300454
rect 407146 300218 407382 300454
rect 406826 299898 407062 300134
rect 407146 299898 407382 300134
rect 406826 264218 407062 264454
rect 407146 264218 407382 264454
rect 406826 263898 407062 264134
rect 407146 263898 407382 264134
rect 406826 228218 407062 228454
rect 407146 228218 407382 228454
rect 406826 227898 407062 228134
rect 407146 227898 407382 228134
rect 406826 192218 407062 192454
rect 407146 192218 407382 192454
rect 406826 191898 407062 192134
rect 407146 191898 407382 192134
rect 406826 156218 407062 156454
rect 407146 156218 407382 156454
rect 406826 155898 407062 156134
rect 407146 155898 407382 156134
rect 406826 120218 407062 120454
rect 407146 120218 407382 120454
rect 406826 119898 407062 120134
rect 407146 119898 407382 120134
rect 406826 84218 407062 84454
rect 407146 84218 407382 84454
rect 406826 83898 407062 84134
rect 407146 83898 407382 84134
rect 406826 48218 407062 48454
rect 407146 48218 407382 48454
rect 406826 47898 407062 48134
rect 407146 47898 407382 48134
rect 406826 12218 407062 12454
rect 407146 12218 407382 12454
rect 406826 11898 407062 12134
rect 407146 11898 407382 12134
rect 406826 -2502 407062 -2266
rect 407146 -2502 407382 -2266
rect 406826 -2822 407062 -2586
rect 407146 -2822 407382 -2586
rect 411326 484718 411562 484954
rect 411646 484718 411882 484954
rect 411326 484398 411562 484634
rect 411646 484398 411882 484634
rect 411326 448718 411562 448954
rect 411646 448718 411882 448954
rect 411326 448398 411562 448634
rect 411646 448398 411882 448634
rect 411326 412718 411562 412954
rect 411646 412718 411882 412954
rect 411326 412398 411562 412634
rect 411646 412398 411882 412634
rect 411326 376718 411562 376954
rect 411646 376718 411882 376954
rect 411326 376398 411562 376634
rect 411646 376398 411882 376634
rect 411326 340718 411562 340954
rect 411646 340718 411882 340954
rect 411326 340398 411562 340634
rect 411646 340398 411882 340634
rect 411326 304718 411562 304954
rect 411646 304718 411882 304954
rect 411326 304398 411562 304634
rect 411646 304398 411882 304634
rect 411326 268718 411562 268954
rect 411646 268718 411882 268954
rect 411326 268398 411562 268634
rect 411646 268398 411882 268634
rect 411326 232718 411562 232954
rect 411646 232718 411882 232954
rect 411326 232398 411562 232634
rect 411646 232398 411882 232634
rect 411326 196718 411562 196954
rect 411646 196718 411882 196954
rect 411326 196398 411562 196634
rect 411646 196398 411882 196634
rect 411326 160718 411562 160954
rect 411646 160718 411882 160954
rect 411326 160398 411562 160634
rect 411646 160398 411882 160634
rect 411326 124718 411562 124954
rect 411646 124718 411882 124954
rect 411326 124398 411562 124634
rect 411646 124398 411882 124634
rect 411326 88718 411562 88954
rect 411646 88718 411882 88954
rect 411326 88398 411562 88634
rect 411646 88398 411882 88634
rect 411326 52718 411562 52954
rect 411646 52718 411882 52954
rect 411326 52398 411562 52634
rect 411646 52398 411882 52634
rect 411326 16718 411562 16954
rect 411646 16718 411882 16954
rect 411326 16398 411562 16634
rect 411646 16398 411882 16634
rect 411326 -3462 411562 -3226
rect 411646 -3462 411882 -3226
rect 411326 -3782 411562 -3546
rect 411646 -3782 411882 -3546
rect 415826 489218 416062 489454
rect 416146 489218 416382 489454
rect 415826 488898 416062 489134
rect 416146 488898 416382 489134
rect 415826 453218 416062 453454
rect 416146 453218 416382 453454
rect 415826 452898 416062 453134
rect 416146 452898 416382 453134
rect 415826 417218 416062 417454
rect 416146 417218 416382 417454
rect 415826 416898 416062 417134
rect 416146 416898 416382 417134
rect 415826 381218 416062 381454
rect 416146 381218 416382 381454
rect 415826 380898 416062 381134
rect 416146 380898 416382 381134
rect 415826 345218 416062 345454
rect 416146 345218 416382 345454
rect 415826 344898 416062 345134
rect 416146 344898 416382 345134
rect 415826 309218 416062 309454
rect 416146 309218 416382 309454
rect 415826 308898 416062 309134
rect 416146 308898 416382 309134
rect 415826 273218 416062 273454
rect 416146 273218 416382 273454
rect 415826 272898 416062 273134
rect 416146 272898 416382 273134
rect 415826 237218 416062 237454
rect 416146 237218 416382 237454
rect 415826 236898 416062 237134
rect 416146 236898 416382 237134
rect 415826 201218 416062 201454
rect 416146 201218 416382 201454
rect 415826 200898 416062 201134
rect 416146 200898 416382 201134
rect 415826 165218 416062 165454
rect 416146 165218 416382 165454
rect 415826 164898 416062 165134
rect 416146 164898 416382 165134
rect 415826 129218 416062 129454
rect 416146 129218 416382 129454
rect 415826 128898 416062 129134
rect 416146 128898 416382 129134
rect 415826 93218 416062 93454
rect 416146 93218 416382 93454
rect 415826 92898 416062 93134
rect 416146 92898 416382 93134
rect 415826 57218 416062 57454
rect 416146 57218 416382 57454
rect 415826 56898 416062 57134
rect 416146 56898 416382 57134
rect 415826 21218 416062 21454
rect 416146 21218 416382 21454
rect 415826 20898 416062 21134
rect 416146 20898 416382 21134
rect 415826 -4422 416062 -4186
rect 416146 -4422 416382 -4186
rect 415826 -4742 416062 -4506
rect 416146 -4742 416382 -4506
rect 420326 493718 420562 493954
rect 420646 493718 420882 493954
rect 420326 493398 420562 493634
rect 420646 493398 420882 493634
rect 420326 457718 420562 457954
rect 420646 457718 420882 457954
rect 420326 457398 420562 457634
rect 420646 457398 420882 457634
rect 420326 421718 420562 421954
rect 420646 421718 420882 421954
rect 420326 421398 420562 421634
rect 420646 421398 420882 421634
rect 420326 385718 420562 385954
rect 420646 385718 420882 385954
rect 420326 385398 420562 385634
rect 420646 385398 420882 385634
rect 420326 349718 420562 349954
rect 420646 349718 420882 349954
rect 420326 349398 420562 349634
rect 420646 349398 420882 349634
rect 420326 313718 420562 313954
rect 420646 313718 420882 313954
rect 420326 313398 420562 313634
rect 420646 313398 420882 313634
rect 420326 277718 420562 277954
rect 420646 277718 420882 277954
rect 420326 277398 420562 277634
rect 420646 277398 420882 277634
rect 420326 241718 420562 241954
rect 420646 241718 420882 241954
rect 420326 241398 420562 241634
rect 420646 241398 420882 241634
rect 420326 205718 420562 205954
rect 420646 205718 420882 205954
rect 420326 205398 420562 205634
rect 420646 205398 420882 205634
rect 420326 169718 420562 169954
rect 420646 169718 420882 169954
rect 420326 169398 420562 169634
rect 420646 169398 420882 169634
rect 420326 133718 420562 133954
rect 420646 133718 420882 133954
rect 420326 133398 420562 133634
rect 420646 133398 420882 133634
rect 420326 97718 420562 97954
rect 420646 97718 420882 97954
rect 420326 97398 420562 97634
rect 420646 97398 420882 97634
rect 420326 61718 420562 61954
rect 420646 61718 420882 61954
rect 420326 61398 420562 61634
rect 420646 61398 420882 61634
rect 420326 25718 420562 25954
rect 420646 25718 420882 25954
rect 420326 25398 420562 25634
rect 420646 25398 420882 25634
rect 420326 -5382 420562 -5146
rect 420646 -5382 420882 -5146
rect 420326 -5702 420562 -5466
rect 420646 -5702 420882 -5466
rect 424826 462218 425062 462454
rect 425146 462218 425382 462454
rect 424826 461898 425062 462134
rect 425146 461898 425382 462134
rect 424826 426218 425062 426454
rect 425146 426218 425382 426454
rect 424826 425898 425062 426134
rect 425146 425898 425382 426134
rect 424826 390218 425062 390454
rect 425146 390218 425382 390454
rect 424826 389898 425062 390134
rect 425146 389898 425382 390134
rect 424826 354218 425062 354454
rect 425146 354218 425382 354454
rect 424826 353898 425062 354134
rect 425146 353898 425382 354134
rect 424826 318218 425062 318454
rect 425146 318218 425382 318454
rect 424826 317898 425062 318134
rect 425146 317898 425382 318134
rect 424826 282218 425062 282454
rect 425146 282218 425382 282454
rect 424826 281898 425062 282134
rect 425146 281898 425382 282134
rect 424826 246218 425062 246454
rect 425146 246218 425382 246454
rect 424826 245898 425062 246134
rect 425146 245898 425382 246134
rect 424826 210218 425062 210454
rect 425146 210218 425382 210454
rect 424826 209898 425062 210134
rect 425146 209898 425382 210134
rect 424826 174218 425062 174454
rect 425146 174218 425382 174454
rect 424826 173898 425062 174134
rect 425146 173898 425382 174134
rect 424826 138218 425062 138454
rect 425146 138218 425382 138454
rect 424826 137898 425062 138134
rect 425146 137898 425382 138134
rect 424826 102218 425062 102454
rect 425146 102218 425382 102454
rect 424826 101898 425062 102134
rect 425146 101898 425382 102134
rect 424826 66218 425062 66454
rect 425146 66218 425382 66454
rect 424826 65898 425062 66134
rect 425146 65898 425382 66134
rect 424826 30218 425062 30454
rect 425146 30218 425382 30454
rect 424826 29898 425062 30134
rect 425146 29898 425382 30134
rect 424826 -6342 425062 -6106
rect 425146 -6342 425382 -6106
rect 424826 -6662 425062 -6426
rect 425146 -6662 425382 -6426
rect 429326 466718 429562 466954
rect 429646 466718 429882 466954
rect 429326 466398 429562 466634
rect 429646 466398 429882 466634
rect 429326 430718 429562 430954
rect 429646 430718 429882 430954
rect 429326 430398 429562 430634
rect 429646 430398 429882 430634
rect 429326 394718 429562 394954
rect 429646 394718 429882 394954
rect 429326 394398 429562 394634
rect 429646 394398 429882 394634
rect 429326 358718 429562 358954
rect 429646 358718 429882 358954
rect 429326 358398 429562 358634
rect 429646 358398 429882 358634
rect 429326 322718 429562 322954
rect 429646 322718 429882 322954
rect 429326 322398 429562 322634
rect 429646 322398 429882 322634
rect 429326 286718 429562 286954
rect 429646 286718 429882 286954
rect 429326 286398 429562 286634
rect 429646 286398 429882 286634
rect 429326 250718 429562 250954
rect 429646 250718 429882 250954
rect 429326 250398 429562 250634
rect 429646 250398 429882 250634
rect 429326 214718 429562 214954
rect 429646 214718 429882 214954
rect 429326 214398 429562 214634
rect 429646 214398 429882 214634
rect 429326 178718 429562 178954
rect 429646 178718 429882 178954
rect 429326 178398 429562 178634
rect 429646 178398 429882 178634
rect 429326 142718 429562 142954
rect 429646 142718 429882 142954
rect 429326 142398 429562 142634
rect 429646 142398 429882 142634
rect 429326 106718 429562 106954
rect 429646 106718 429882 106954
rect 429326 106398 429562 106634
rect 429646 106398 429882 106634
rect 429326 70718 429562 70954
rect 429646 70718 429882 70954
rect 429326 70398 429562 70634
rect 429646 70398 429882 70634
rect 429326 34718 429562 34954
rect 429646 34718 429882 34954
rect 429326 34398 429562 34634
rect 429646 34398 429882 34634
rect 429326 -7302 429562 -7066
rect 429646 -7302 429882 -7066
rect 429326 -7622 429562 -7386
rect 429646 -7622 429882 -7386
rect 433826 471218 434062 471454
rect 434146 471218 434382 471454
rect 433826 470898 434062 471134
rect 434146 470898 434382 471134
rect 433826 435218 434062 435454
rect 434146 435218 434382 435454
rect 433826 434898 434062 435134
rect 434146 434898 434382 435134
rect 433826 399218 434062 399454
rect 434146 399218 434382 399454
rect 433826 398898 434062 399134
rect 434146 398898 434382 399134
rect 433826 363218 434062 363454
rect 434146 363218 434382 363454
rect 433826 362898 434062 363134
rect 434146 362898 434382 363134
rect 433826 327218 434062 327454
rect 434146 327218 434382 327454
rect 433826 326898 434062 327134
rect 434146 326898 434382 327134
rect 433826 291218 434062 291454
rect 434146 291218 434382 291454
rect 433826 290898 434062 291134
rect 434146 290898 434382 291134
rect 433826 255218 434062 255454
rect 434146 255218 434382 255454
rect 433826 254898 434062 255134
rect 434146 254898 434382 255134
rect 433826 219218 434062 219454
rect 434146 219218 434382 219454
rect 433826 218898 434062 219134
rect 434146 218898 434382 219134
rect 433826 183218 434062 183454
rect 434146 183218 434382 183454
rect 433826 182898 434062 183134
rect 434146 182898 434382 183134
rect 433826 147218 434062 147454
rect 434146 147218 434382 147454
rect 433826 146898 434062 147134
rect 434146 146898 434382 147134
rect 433826 111218 434062 111454
rect 434146 111218 434382 111454
rect 433826 110898 434062 111134
rect 434146 110898 434382 111134
rect 433826 75218 434062 75454
rect 434146 75218 434382 75454
rect 433826 74898 434062 75134
rect 434146 74898 434382 75134
rect 433826 39218 434062 39454
rect 434146 39218 434382 39454
rect 433826 38898 434062 39134
rect 434146 38898 434382 39134
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 438326 475718 438562 475954
rect 438646 475718 438882 475954
rect 438326 475398 438562 475634
rect 438646 475398 438882 475634
rect 438326 439718 438562 439954
rect 438646 439718 438882 439954
rect 438326 439398 438562 439634
rect 438646 439398 438882 439634
rect 438326 403718 438562 403954
rect 438646 403718 438882 403954
rect 438326 403398 438562 403634
rect 438646 403398 438882 403634
rect 438326 367718 438562 367954
rect 438646 367718 438882 367954
rect 438326 367398 438562 367634
rect 438646 367398 438882 367634
rect 438326 331718 438562 331954
rect 438646 331718 438882 331954
rect 438326 331398 438562 331634
rect 438646 331398 438882 331634
rect 438326 295718 438562 295954
rect 438646 295718 438882 295954
rect 438326 295398 438562 295634
rect 438646 295398 438882 295634
rect 438326 259718 438562 259954
rect 438646 259718 438882 259954
rect 438326 259398 438562 259634
rect 438646 259398 438882 259634
rect 438326 223718 438562 223954
rect 438646 223718 438882 223954
rect 438326 223398 438562 223634
rect 438646 223398 438882 223634
rect 438326 187718 438562 187954
rect 438646 187718 438882 187954
rect 438326 187398 438562 187634
rect 438646 187398 438882 187634
rect 438326 151718 438562 151954
rect 438646 151718 438882 151954
rect 438326 151398 438562 151634
rect 438646 151398 438882 151634
rect 438326 115718 438562 115954
rect 438646 115718 438882 115954
rect 438326 115398 438562 115634
rect 438646 115398 438882 115634
rect 438326 79718 438562 79954
rect 438646 79718 438882 79954
rect 438326 79398 438562 79634
rect 438646 79398 438882 79634
rect 438326 43718 438562 43954
rect 438646 43718 438882 43954
rect 438326 43398 438562 43634
rect 438646 43398 438882 43634
rect 438326 7718 438562 7954
rect 438646 7718 438882 7954
rect 438326 7398 438562 7634
rect 438646 7398 438882 7634
rect 438326 -1542 438562 -1306
rect 438646 -1542 438882 -1306
rect 438326 -1862 438562 -1626
rect 438646 -1862 438882 -1626
rect 442826 480218 443062 480454
rect 443146 480218 443382 480454
rect 442826 479898 443062 480134
rect 443146 479898 443382 480134
rect 442826 444218 443062 444454
rect 443146 444218 443382 444454
rect 442826 443898 443062 444134
rect 443146 443898 443382 444134
rect 442826 408218 443062 408454
rect 443146 408218 443382 408454
rect 442826 407898 443062 408134
rect 443146 407898 443382 408134
rect 442826 372218 443062 372454
rect 443146 372218 443382 372454
rect 442826 371898 443062 372134
rect 443146 371898 443382 372134
rect 442826 336218 443062 336454
rect 443146 336218 443382 336454
rect 442826 335898 443062 336134
rect 443146 335898 443382 336134
rect 442826 300218 443062 300454
rect 443146 300218 443382 300454
rect 442826 299898 443062 300134
rect 443146 299898 443382 300134
rect 442826 264218 443062 264454
rect 443146 264218 443382 264454
rect 442826 263898 443062 264134
rect 443146 263898 443382 264134
rect 442826 228218 443062 228454
rect 443146 228218 443382 228454
rect 442826 227898 443062 228134
rect 443146 227898 443382 228134
rect 442826 192218 443062 192454
rect 443146 192218 443382 192454
rect 442826 191898 443062 192134
rect 443146 191898 443382 192134
rect 442826 156218 443062 156454
rect 443146 156218 443382 156454
rect 442826 155898 443062 156134
rect 443146 155898 443382 156134
rect 442826 120218 443062 120454
rect 443146 120218 443382 120454
rect 442826 119898 443062 120134
rect 443146 119898 443382 120134
rect 442826 84218 443062 84454
rect 443146 84218 443382 84454
rect 442826 83898 443062 84134
rect 443146 83898 443382 84134
rect 442826 48218 443062 48454
rect 443146 48218 443382 48454
rect 442826 47898 443062 48134
rect 443146 47898 443382 48134
rect 442826 12218 443062 12454
rect 443146 12218 443382 12454
rect 442826 11898 443062 12134
rect 443146 11898 443382 12134
rect 442826 -2502 443062 -2266
rect 443146 -2502 443382 -2266
rect 442826 -2822 443062 -2586
rect 443146 -2822 443382 -2586
rect 447326 484718 447562 484954
rect 447646 484718 447882 484954
rect 447326 484398 447562 484634
rect 447646 484398 447882 484634
rect 447326 448718 447562 448954
rect 447646 448718 447882 448954
rect 447326 448398 447562 448634
rect 447646 448398 447882 448634
rect 447326 412718 447562 412954
rect 447646 412718 447882 412954
rect 447326 412398 447562 412634
rect 447646 412398 447882 412634
rect 447326 376718 447562 376954
rect 447646 376718 447882 376954
rect 447326 376398 447562 376634
rect 447646 376398 447882 376634
rect 447326 340718 447562 340954
rect 447646 340718 447882 340954
rect 447326 340398 447562 340634
rect 447646 340398 447882 340634
rect 447326 304718 447562 304954
rect 447646 304718 447882 304954
rect 447326 304398 447562 304634
rect 447646 304398 447882 304634
rect 447326 268718 447562 268954
rect 447646 268718 447882 268954
rect 447326 268398 447562 268634
rect 447646 268398 447882 268634
rect 447326 232718 447562 232954
rect 447646 232718 447882 232954
rect 447326 232398 447562 232634
rect 447646 232398 447882 232634
rect 447326 196718 447562 196954
rect 447646 196718 447882 196954
rect 447326 196398 447562 196634
rect 447646 196398 447882 196634
rect 447326 160718 447562 160954
rect 447646 160718 447882 160954
rect 447326 160398 447562 160634
rect 447646 160398 447882 160634
rect 447326 124718 447562 124954
rect 447646 124718 447882 124954
rect 447326 124398 447562 124634
rect 447646 124398 447882 124634
rect 447326 88718 447562 88954
rect 447646 88718 447882 88954
rect 447326 88398 447562 88634
rect 447646 88398 447882 88634
rect 447326 52718 447562 52954
rect 447646 52718 447882 52954
rect 447326 52398 447562 52634
rect 447646 52398 447882 52634
rect 447326 16718 447562 16954
rect 447646 16718 447882 16954
rect 447326 16398 447562 16634
rect 447646 16398 447882 16634
rect 447326 -3462 447562 -3226
rect 447646 -3462 447882 -3226
rect 447326 -3782 447562 -3546
rect 447646 -3782 447882 -3546
rect 451826 489218 452062 489454
rect 452146 489218 452382 489454
rect 451826 488898 452062 489134
rect 452146 488898 452382 489134
rect 451826 453218 452062 453454
rect 452146 453218 452382 453454
rect 451826 452898 452062 453134
rect 452146 452898 452382 453134
rect 451826 417218 452062 417454
rect 452146 417218 452382 417454
rect 451826 416898 452062 417134
rect 452146 416898 452382 417134
rect 451826 381218 452062 381454
rect 452146 381218 452382 381454
rect 451826 380898 452062 381134
rect 452146 380898 452382 381134
rect 451826 345218 452062 345454
rect 452146 345218 452382 345454
rect 451826 344898 452062 345134
rect 452146 344898 452382 345134
rect 451826 309218 452062 309454
rect 452146 309218 452382 309454
rect 451826 308898 452062 309134
rect 452146 308898 452382 309134
rect 451826 273218 452062 273454
rect 452146 273218 452382 273454
rect 451826 272898 452062 273134
rect 452146 272898 452382 273134
rect 451826 237218 452062 237454
rect 452146 237218 452382 237454
rect 451826 236898 452062 237134
rect 452146 236898 452382 237134
rect 451826 201218 452062 201454
rect 452146 201218 452382 201454
rect 451826 200898 452062 201134
rect 452146 200898 452382 201134
rect 451826 165218 452062 165454
rect 452146 165218 452382 165454
rect 451826 164898 452062 165134
rect 452146 164898 452382 165134
rect 451826 129218 452062 129454
rect 452146 129218 452382 129454
rect 451826 128898 452062 129134
rect 452146 128898 452382 129134
rect 451826 93218 452062 93454
rect 452146 93218 452382 93454
rect 451826 92898 452062 93134
rect 452146 92898 452382 93134
rect 451826 57218 452062 57454
rect 452146 57218 452382 57454
rect 451826 56898 452062 57134
rect 452146 56898 452382 57134
rect 451826 21218 452062 21454
rect 452146 21218 452382 21454
rect 451826 20898 452062 21134
rect 452146 20898 452382 21134
rect 451826 -4422 452062 -4186
rect 452146 -4422 452382 -4186
rect 451826 -4742 452062 -4506
rect 452146 -4742 452382 -4506
rect 456326 493718 456562 493954
rect 456646 493718 456882 493954
rect 456326 493398 456562 493634
rect 456646 493398 456882 493634
rect 456326 457718 456562 457954
rect 456646 457718 456882 457954
rect 456326 457398 456562 457634
rect 456646 457398 456882 457634
rect 456326 421718 456562 421954
rect 456646 421718 456882 421954
rect 456326 421398 456562 421634
rect 456646 421398 456882 421634
rect 456326 385718 456562 385954
rect 456646 385718 456882 385954
rect 456326 385398 456562 385634
rect 456646 385398 456882 385634
rect 456326 349718 456562 349954
rect 456646 349718 456882 349954
rect 456326 349398 456562 349634
rect 456646 349398 456882 349634
rect 456326 313718 456562 313954
rect 456646 313718 456882 313954
rect 456326 313398 456562 313634
rect 456646 313398 456882 313634
rect 456326 277718 456562 277954
rect 456646 277718 456882 277954
rect 456326 277398 456562 277634
rect 456646 277398 456882 277634
rect 456326 241718 456562 241954
rect 456646 241718 456882 241954
rect 456326 241398 456562 241634
rect 456646 241398 456882 241634
rect 456326 205718 456562 205954
rect 456646 205718 456882 205954
rect 456326 205398 456562 205634
rect 456646 205398 456882 205634
rect 456326 169718 456562 169954
rect 456646 169718 456882 169954
rect 456326 169398 456562 169634
rect 456646 169398 456882 169634
rect 456326 133718 456562 133954
rect 456646 133718 456882 133954
rect 456326 133398 456562 133634
rect 456646 133398 456882 133634
rect 456326 97718 456562 97954
rect 456646 97718 456882 97954
rect 456326 97398 456562 97634
rect 456646 97398 456882 97634
rect 456326 61718 456562 61954
rect 456646 61718 456882 61954
rect 456326 61398 456562 61634
rect 456646 61398 456882 61634
rect 456326 25718 456562 25954
rect 456646 25718 456882 25954
rect 456326 25398 456562 25634
rect 456646 25398 456882 25634
rect 456326 -5382 456562 -5146
rect 456646 -5382 456882 -5146
rect 456326 -5702 456562 -5466
rect 456646 -5702 456882 -5466
rect 460826 462218 461062 462454
rect 461146 462218 461382 462454
rect 460826 461898 461062 462134
rect 461146 461898 461382 462134
rect 460826 426218 461062 426454
rect 461146 426218 461382 426454
rect 460826 425898 461062 426134
rect 461146 425898 461382 426134
rect 460826 390218 461062 390454
rect 461146 390218 461382 390454
rect 460826 389898 461062 390134
rect 461146 389898 461382 390134
rect 460826 354218 461062 354454
rect 461146 354218 461382 354454
rect 460826 353898 461062 354134
rect 461146 353898 461382 354134
rect 460826 318218 461062 318454
rect 461146 318218 461382 318454
rect 460826 317898 461062 318134
rect 461146 317898 461382 318134
rect 460826 282218 461062 282454
rect 461146 282218 461382 282454
rect 460826 281898 461062 282134
rect 461146 281898 461382 282134
rect 460826 246218 461062 246454
rect 461146 246218 461382 246454
rect 460826 245898 461062 246134
rect 461146 245898 461382 246134
rect 460826 210218 461062 210454
rect 461146 210218 461382 210454
rect 460826 209898 461062 210134
rect 461146 209898 461382 210134
rect 460826 174218 461062 174454
rect 461146 174218 461382 174454
rect 460826 173898 461062 174134
rect 461146 173898 461382 174134
rect 460826 138218 461062 138454
rect 461146 138218 461382 138454
rect 460826 137898 461062 138134
rect 461146 137898 461382 138134
rect 460826 102218 461062 102454
rect 461146 102218 461382 102454
rect 460826 101898 461062 102134
rect 461146 101898 461382 102134
rect 460826 66218 461062 66454
rect 461146 66218 461382 66454
rect 460826 65898 461062 66134
rect 461146 65898 461382 66134
rect 460826 30218 461062 30454
rect 461146 30218 461382 30454
rect 460826 29898 461062 30134
rect 461146 29898 461382 30134
rect 460826 -6342 461062 -6106
rect 461146 -6342 461382 -6106
rect 460826 -6662 461062 -6426
rect 461146 -6662 461382 -6426
rect 465326 466718 465562 466954
rect 465646 466718 465882 466954
rect 465326 466398 465562 466634
rect 465646 466398 465882 466634
rect 465326 430718 465562 430954
rect 465646 430718 465882 430954
rect 465326 430398 465562 430634
rect 465646 430398 465882 430634
rect 465326 394718 465562 394954
rect 465646 394718 465882 394954
rect 465326 394398 465562 394634
rect 465646 394398 465882 394634
rect 465326 358718 465562 358954
rect 465646 358718 465882 358954
rect 465326 358398 465562 358634
rect 465646 358398 465882 358634
rect 465326 322718 465562 322954
rect 465646 322718 465882 322954
rect 465326 322398 465562 322634
rect 465646 322398 465882 322634
rect 465326 286718 465562 286954
rect 465646 286718 465882 286954
rect 465326 286398 465562 286634
rect 465646 286398 465882 286634
rect 465326 250718 465562 250954
rect 465646 250718 465882 250954
rect 465326 250398 465562 250634
rect 465646 250398 465882 250634
rect 465326 214718 465562 214954
rect 465646 214718 465882 214954
rect 465326 214398 465562 214634
rect 465646 214398 465882 214634
rect 465326 178718 465562 178954
rect 465646 178718 465882 178954
rect 465326 178398 465562 178634
rect 465646 178398 465882 178634
rect 465326 142718 465562 142954
rect 465646 142718 465882 142954
rect 465326 142398 465562 142634
rect 465646 142398 465882 142634
rect 465326 106718 465562 106954
rect 465646 106718 465882 106954
rect 465326 106398 465562 106634
rect 465646 106398 465882 106634
rect 465326 70718 465562 70954
rect 465646 70718 465882 70954
rect 465326 70398 465562 70634
rect 465646 70398 465882 70634
rect 465326 34718 465562 34954
rect 465646 34718 465882 34954
rect 465326 34398 465562 34634
rect 465646 34398 465882 34634
rect 465326 -7302 465562 -7066
rect 465646 -7302 465882 -7066
rect 465326 -7622 465562 -7386
rect 465646 -7622 465882 -7386
rect 469826 471218 470062 471454
rect 470146 471218 470382 471454
rect 469826 470898 470062 471134
rect 470146 470898 470382 471134
rect 469826 435218 470062 435454
rect 470146 435218 470382 435454
rect 469826 434898 470062 435134
rect 470146 434898 470382 435134
rect 469826 399218 470062 399454
rect 470146 399218 470382 399454
rect 469826 398898 470062 399134
rect 470146 398898 470382 399134
rect 469826 363218 470062 363454
rect 470146 363218 470382 363454
rect 469826 362898 470062 363134
rect 470146 362898 470382 363134
rect 469826 327218 470062 327454
rect 470146 327218 470382 327454
rect 469826 326898 470062 327134
rect 470146 326898 470382 327134
rect 469826 291218 470062 291454
rect 470146 291218 470382 291454
rect 469826 290898 470062 291134
rect 470146 290898 470382 291134
rect 469826 255218 470062 255454
rect 470146 255218 470382 255454
rect 469826 254898 470062 255134
rect 470146 254898 470382 255134
rect 469826 219218 470062 219454
rect 470146 219218 470382 219454
rect 469826 218898 470062 219134
rect 470146 218898 470382 219134
rect 469826 183218 470062 183454
rect 470146 183218 470382 183454
rect 469826 182898 470062 183134
rect 470146 182898 470382 183134
rect 469826 147218 470062 147454
rect 470146 147218 470382 147454
rect 469826 146898 470062 147134
rect 470146 146898 470382 147134
rect 469826 111218 470062 111454
rect 470146 111218 470382 111454
rect 469826 110898 470062 111134
rect 470146 110898 470382 111134
rect 469826 75218 470062 75454
rect 470146 75218 470382 75454
rect 469826 74898 470062 75134
rect 470146 74898 470382 75134
rect 469826 39218 470062 39454
rect 470146 39218 470382 39454
rect 469826 38898 470062 39134
rect 470146 38898 470382 39134
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 474326 475718 474562 475954
rect 474646 475718 474882 475954
rect 474326 475398 474562 475634
rect 474646 475398 474882 475634
rect 474326 439718 474562 439954
rect 474646 439718 474882 439954
rect 474326 439398 474562 439634
rect 474646 439398 474882 439634
rect 474326 403718 474562 403954
rect 474646 403718 474882 403954
rect 474326 403398 474562 403634
rect 474646 403398 474882 403634
rect 474326 367718 474562 367954
rect 474646 367718 474882 367954
rect 474326 367398 474562 367634
rect 474646 367398 474882 367634
rect 474326 331718 474562 331954
rect 474646 331718 474882 331954
rect 474326 331398 474562 331634
rect 474646 331398 474882 331634
rect 474326 295718 474562 295954
rect 474646 295718 474882 295954
rect 474326 295398 474562 295634
rect 474646 295398 474882 295634
rect 474326 259718 474562 259954
rect 474646 259718 474882 259954
rect 474326 259398 474562 259634
rect 474646 259398 474882 259634
rect 474326 223718 474562 223954
rect 474646 223718 474882 223954
rect 474326 223398 474562 223634
rect 474646 223398 474882 223634
rect 474326 187718 474562 187954
rect 474646 187718 474882 187954
rect 474326 187398 474562 187634
rect 474646 187398 474882 187634
rect 474326 151718 474562 151954
rect 474646 151718 474882 151954
rect 474326 151398 474562 151634
rect 474646 151398 474882 151634
rect 474326 115718 474562 115954
rect 474646 115718 474882 115954
rect 474326 115398 474562 115634
rect 474646 115398 474882 115634
rect 474326 79718 474562 79954
rect 474646 79718 474882 79954
rect 474326 79398 474562 79634
rect 474646 79398 474882 79634
rect 474326 43718 474562 43954
rect 474646 43718 474882 43954
rect 474326 43398 474562 43634
rect 474646 43398 474882 43634
rect 474326 7718 474562 7954
rect 474646 7718 474882 7954
rect 474326 7398 474562 7634
rect 474646 7398 474882 7634
rect 474326 -1542 474562 -1306
rect 474646 -1542 474882 -1306
rect 474326 -1862 474562 -1626
rect 474646 -1862 474882 -1626
rect 478826 706522 479062 706758
rect 479146 706522 479382 706758
rect 478826 706202 479062 706438
rect 479146 706202 479382 706438
rect 478826 696218 479062 696454
rect 479146 696218 479382 696454
rect 478826 695898 479062 696134
rect 479146 695898 479382 696134
rect 478826 660218 479062 660454
rect 479146 660218 479382 660454
rect 478826 659898 479062 660134
rect 479146 659898 479382 660134
rect 478826 624218 479062 624454
rect 479146 624218 479382 624454
rect 478826 623898 479062 624134
rect 479146 623898 479382 624134
rect 478826 588218 479062 588454
rect 479146 588218 479382 588454
rect 478826 587898 479062 588134
rect 479146 587898 479382 588134
rect 478826 552218 479062 552454
rect 479146 552218 479382 552454
rect 478826 551898 479062 552134
rect 479146 551898 479382 552134
rect 478826 516218 479062 516454
rect 479146 516218 479382 516454
rect 478826 515898 479062 516134
rect 479146 515898 479382 516134
rect 478826 480218 479062 480454
rect 479146 480218 479382 480454
rect 478826 479898 479062 480134
rect 479146 479898 479382 480134
rect 478826 444218 479062 444454
rect 479146 444218 479382 444454
rect 478826 443898 479062 444134
rect 479146 443898 479382 444134
rect 478826 408218 479062 408454
rect 479146 408218 479382 408454
rect 478826 407898 479062 408134
rect 479146 407898 479382 408134
rect 478826 372218 479062 372454
rect 479146 372218 479382 372454
rect 478826 371898 479062 372134
rect 479146 371898 479382 372134
rect 478826 336218 479062 336454
rect 479146 336218 479382 336454
rect 478826 335898 479062 336134
rect 479146 335898 479382 336134
rect 478826 300218 479062 300454
rect 479146 300218 479382 300454
rect 478826 299898 479062 300134
rect 479146 299898 479382 300134
rect 478826 264218 479062 264454
rect 479146 264218 479382 264454
rect 478826 263898 479062 264134
rect 479146 263898 479382 264134
rect 478826 228218 479062 228454
rect 479146 228218 479382 228454
rect 478826 227898 479062 228134
rect 479146 227898 479382 228134
rect 478826 192218 479062 192454
rect 479146 192218 479382 192454
rect 478826 191898 479062 192134
rect 479146 191898 479382 192134
rect 478826 156218 479062 156454
rect 479146 156218 479382 156454
rect 478826 155898 479062 156134
rect 479146 155898 479382 156134
rect 478826 120218 479062 120454
rect 479146 120218 479382 120454
rect 478826 119898 479062 120134
rect 479146 119898 479382 120134
rect 478826 84218 479062 84454
rect 479146 84218 479382 84454
rect 478826 83898 479062 84134
rect 479146 83898 479382 84134
rect 478826 48218 479062 48454
rect 479146 48218 479382 48454
rect 478826 47898 479062 48134
rect 479146 47898 479382 48134
rect 478826 12218 479062 12454
rect 479146 12218 479382 12454
rect 478826 11898 479062 12134
rect 479146 11898 479382 12134
rect 478826 -2502 479062 -2266
rect 479146 -2502 479382 -2266
rect 478826 -2822 479062 -2586
rect 479146 -2822 479382 -2586
rect 483326 707482 483562 707718
rect 483646 707482 483882 707718
rect 483326 707162 483562 707398
rect 483646 707162 483882 707398
rect 483326 700718 483562 700954
rect 483646 700718 483882 700954
rect 483326 700398 483562 700634
rect 483646 700398 483882 700634
rect 483326 664718 483562 664954
rect 483646 664718 483882 664954
rect 483326 664398 483562 664634
rect 483646 664398 483882 664634
rect 483326 628718 483562 628954
rect 483646 628718 483882 628954
rect 483326 628398 483562 628634
rect 483646 628398 483882 628634
rect 483326 592718 483562 592954
rect 483646 592718 483882 592954
rect 483326 592398 483562 592634
rect 483646 592398 483882 592634
rect 483326 556718 483562 556954
rect 483646 556718 483882 556954
rect 483326 556398 483562 556634
rect 483646 556398 483882 556634
rect 483326 520718 483562 520954
rect 483646 520718 483882 520954
rect 483326 520398 483562 520634
rect 483646 520398 483882 520634
rect 483326 484718 483562 484954
rect 483646 484718 483882 484954
rect 483326 484398 483562 484634
rect 483646 484398 483882 484634
rect 483326 448718 483562 448954
rect 483646 448718 483882 448954
rect 483326 448398 483562 448634
rect 483646 448398 483882 448634
rect 483326 412718 483562 412954
rect 483646 412718 483882 412954
rect 483326 412398 483562 412634
rect 483646 412398 483882 412634
rect 483326 376718 483562 376954
rect 483646 376718 483882 376954
rect 483326 376398 483562 376634
rect 483646 376398 483882 376634
rect 483326 340718 483562 340954
rect 483646 340718 483882 340954
rect 483326 340398 483562 340634
rect 483646 340398 483882 340634
rect 483326 304718 483562 304954
rect 483646 304718 483882 304954
rect 483326 304398 483562 304634
rect 483646 304398 483882 304634
rect 483326 268718 483562 268954
rect 483646 268718 483882 268954
rect 483326 268398 483562 268634
rect 483646 268398 483882 268634
rect 483326 232718 483562 232954
rect 483646 232718 483882 232954
rect 483326 232398 483562 232634
rect 483646 232398 483882 232634
rect 483326 196718 483562 196954
rect 483646 196718 483882 196954
rect 483326 196398 483562 196634
rect 483646 196398 483882 196634
rect 483326 160718 483562 160954
rect 483646 160718 483882 160954
rect 483326 160398 483562 160634
rect 483646 160398 483882 160634
rect 483326 124718 483562 124954
rect 483646 124718 483882 124954
rect 483326 124398 483562 124634
rect 483646 124398 483882 124634
rect 483326 88718 483562 88954
rect 483646 88718 483882 88954
rect 483326 88398 483562 88634
rect 483646 88398 483882 88634
rect 483326 52718 483562 52954
rect 483646 52718 483882 52954
rect 483326 52398 483562 52634
rect 483646 52398 483882 52634
rect 483326 16718 483562 16954
rect 483646 16718 483882 16954
rect 483326 16398 483562 16634
rect 483646 16398 483882 16634
rect 483326 -3462 483562 -3226
rect 483646 -3462 483882 -3226
rect 483326 -3782 483562 -3546
rect 483646 -3782 483882 -3546
rect 487826 708442 488062 708678
rect 488146 708442 488382 708678
rect 487826 708122 488062 708358
rect 488146 708122 488382 708358
rect 487826 669218 488062 669454
rect 488146 669218 488382 669454
rect 487826 668898 488062 669134
rect 488146 668898 488382 669134
rect 487826 633218 488062 633454
rect 488146 633218 488382 633454
rect 487826 632898 488062 633134
rect 488146 632898 488382 633134
rect 487826 597218 488062 597454
rect 488146 597218 488382 597454
rect 487826 596898 488062 597134
rect 488146 596898 488382 597134
rect 487826 561218 488062 561454
rect 488146 561218 488382 561454
rect 487826 560898 488062 561134
rect 488146 560898 488382 561134
rect 487826 525218 488062 525454
rect 488146 525218 488382 525454
rect 487826 524898 488062 525134
rect 488146 524898 488382 525134
rect 487826 489218 488062 489454
rect 488146 489218 488382 489454
rect 487826 488898 488062 489134
rect 488146 488898 488382 489134
rect 487826 453218 488062 453454
rect 488146 453218 488382 453454
rect 487826 452898 488062 453134
rect 488146 452898 488382 453134
rect 487826 417218 488062 417454
rect 488146 417218 488382 417454
rect 487826 416898 488062 417134
rect 488146 416898 488382 417134
rect 487826 381218 488062 381454
rect 488146 381218 488382 381454
rect 487826 380898 488062 381134
rect 488146 380898 488382 381134
rect 487826 345218 488062 345454
rect 488146 345218 488382 345454
rect 487826 344898 488062 345134
rect 488146 344898 488382 345134
rect 487826 309218 488062 309454
rect 488146 309218 488382 309454
rect 487826 308898 488062 309134
rect 488146 308898 488382 309134
rect 487826 273218 488062 273454
rect 488146 273218 488382 273454
rect 487826 272898 488062 273134
rect 488146 272898 488382 273134
rect 487826 237218 488062 237454
rect 488146 237218 488382 237454
rect 487826 236898 488062 237134
rect 488146 236898 488382 237134
rect 487826 201218 488062 201454
rect 488146 201218 488382 201454
rect 487826 200898 488062 201134
rect 488146 200898 488382 201134
rect 487826 165218 488062 165454
rect 488146 165218 488382 165454
rect 487826 164898 488062 165134
rect 488146 164898 488382 165134
rect 487826 129218 488062 129454
rect 488146 129218 488382 129454
rect 487826 128898 488062 129134
rect 488146 128898 488382 129134
rect 487826 93218 488062 93454
rect 488146 93218 488382 93454
rect 487826 92898 488062 93134
rect 488146 92898 488382 93134
rect 487826 57218 488062 57454
rect 488146 57218 488382 57454
rect 487826 56898 488062 57134
rect 488146 56898 488382 57134
rect 487826 21218 488062 21454
rect 488146 21218 488382 21454
rect 487826 20898 488062 21134
rect 488146 20898 488382 21134
rect 487826 -4422 488062 -4186
rect 488146 -4422 488382 -4186
rect 487826 -4742 488062 -4506
rect 488146 -4742 488382 -4506
rect 492326 709402 492562 709638
rect 492646 709402 492882 709638
rect 492326 709082 492562 709318
rect 492646 709082 492882 709318
rect 492326 673718 492562 673954
rect 492646 673718 492882 673954
rect 492326 673398 492562 673634
rect 492646 673398 492882 673634
rect 492326 637718 492562 637954
rect 492646 637718 492882 637954
rect 492326 637398 492562 637634
rect 492646 637398 492882 637634
rect 492326 601718 492562 601954
rect 492646 601718 492882 601954
rect 492326 601398 492562 601634
rect 492646 601398 492882 601634
rect 492326 565718 492562 565954
rect 492646 565718 492882 565954
rect 492326 565398 492562 565634
rect 492646 565398 492882 565634
rect 492326 529718 492562 529954
rect 492646 529718 492882 529954
rect 492326 529398 492562 529634
rect 492646 529398 492882 529634
rect 492326 493718 492562 493954
rect 492646 493718 492882 493954
rect 492326 493398 492562 493634
rect 492646 493398 492882 493634
rect 492326 457718 492562 457954
rect 492646 457718 492882 457954
rect 492326 457398 492562 457634
rect 492646 457398 492882 457634
rect 492326 421718 492562 421954
rect 492646 421718 492882 421954
rect 492326 421398 492562 421634
rect 492646 421398 492882 421634
rect 492326 385718 492562 385954
rect 492646 385718 492882 385954
rect 492326 385398 492562 385634
rect 492646 385398 492882 385634
rect 492326 349718 492562 349954
rect 492646 349718 492882 349954
rect 492326 349398 492562 349634
rect 492646 349398 492882 349634
rect 492326 313718 492562 313954
rect 492646 313718 492882 313954
rect 492326 313398 492562 313634
rect 492646 313398 492882 313634
rect 492326 277718 492562 277954
rect 492646 277718 492882 277954
rect 492326 277398 492562 277634
rect 492646 277398 492882 277634
rect 492326 241718 492562 241954
rect 492646 241718 492882 241954
rect 492326 241398 492562 241634
rect 492646 241398 492882 241634
rect 492326 205718 492562 205954
rect 492646 205718 492882 205954
rect 492326 205398 492562 205634
rect 492646 205398 492882 205634
rect 492326 169718 492562 169954
rect 492646 169718 492882 169954
rect 492326 169398 492562 169634
rect 492646 169398 492882 169634
rect 492326 133718 492562 133954
rect 492646 133718 492882 133954
rect 492326 133398 492562 133634
rect 492646 133398 492882 133634
rect 492326 97718 492562 97954
rect 492646 97718 492882 97954
rect 492326 97398 492562 97634
rect 492646 97398 492882 97634
rect 492326 61718 492562 61954
rect 492646 61718 492882 61954
rect 492326 61398 492562 61634
rect 492646 61398 492882 61634
rect 492326 25718 492562 25954
rect 492646 25718 492882 25954
rect 492326 25398 492562 25634
rect 492646 25398 492882 25634
rect 492326 -5382 492562 -5146
rect 492646 -5382 492882 -5146
rect 492326 -5702 492562 -5466
rect 492646 -5702 492882 -5466
rect 496826 710362 497062 710598
rect 497146 710362 497382 710598
rect 496826 710042 497062 710278
rect 497146 710042 497382 710278
rect 496826 678218 497062 678454
rect 497146 678218 497382 678454
rect 496826 677898 497062 678134
rect 497146 677898 497382 678134
rect 496826 642218 497062 642454
rect 497146 642218 497382 642454
rect 496826 641898 497062 642134
rect 497146 641898 497382 642134
rect 496826 606218 497062 606454
rect 497146 606218 497382 606454
rect 496826 605898 497062 606134
rect 497146 605898 497382 606134
rect 496826 570218 497062 570454
rect 497146 570218 497382 570454
rect 496826 569898 497062 570134
rect 497146 569898 497382 570134
rect 496826 534218 497062 534454
rect 497146 534218 497382 534454
rect 496826 533898 497062 534134
rect 497146 533898 497382 534134
rect 496826 498218 497062 498454
rect 497146 498218 497382 498454
rect 496826 497898 497062 498134
rect 497146 497898 497382 498134
rect 496826 462218 497062 462454
rect 497146 462218 497382 462454
rect 496826 461898 497062 462134
rect 497146 461898 497382 462134
rect 496826 426218 497062 426454
rect 497146 426218 497382 426454
rect 496826 425898 497062 426134
rect 497146 425898 497382 426134
rect 496826 390218 497062 390454
rect 497146 390218 497382 390454
rect 496826 389898 497062 390134
rect 497146 389898 497382 390134
rect 496826 354218 497062 354454
rect 497146 354218 497382 354454
rect 496826 353898 497062 354134
rect 497146 353898 497382 354134
rect 496826 318218 497062 318454
rect 497146 318218 497382 318454
rect 496826 317898 497062 318134
rect 497146 317898 497382 318134
rect 496826 282218 497062 282454
rect 497146 282218 497382 282454
rect 496826 281898 497062 282134
rect 497146 281898 497382 282134
rect 496826 246218 497062 246454
rect 497146 246218 497382 246454
rect 496826 245898 497062 246134
rect 497146 245898 497382 246134
rect 496826 210218 497062 210454
rect 497146 210218 497382 210454
rect 496826 209898 497062 210134
rect 497146 209898 497382 210134
rect 496826 174218 497062 174454
rect 497146 174218 497382 174454
rect 496826 173898 497062 174134
rect 497146 173898 497382 174134
rect 496826 138218 497062 138454
rect 497146 138218 497382 138454
rect 496826 137898 497062 138134
rect 497146 137898 497382 138134
rect 496826 102218 497062 102454
rect 497146 102218 497382 102454
rect 496826 101898 497062 102134
rect 497146 101898 497382 102134
rect 496826 66218 497062 66454
rect 497146 66218 497382 66454
rect 496826 65898 497062 66134
rect 497146 65898 497382 66134
rect 496826 30218 497062 30454
rect 497146 30218 497382 30454
rect 496826 29898 497062 30134
rect 497146 29898 497382 30134
rect 496826 -6342 497062 -6106
rect 497146 -6342 497382 -6106
rect 496826 -6662 497062 -6426
rect 497146 -6662 497382 -6426
rect 501326 711322 501562 711558
rect 501646 711322 501882 711558
rect 501326 711002 501562 711238
rect 501646 711002 501882 711238
rect 501326 682718 501562 682954
rect 501646 682718 501882 682954
rect 501326 682398 501562 682634
rect 501646 682398 501882 682634
rect 501326 646718 501562 646954
rect 501646 646718 501882 646954
rect 501326 646398 501562 646634
rect 501646 646398 501882 646634
rect 501326 610718 501562 610954
rect 501646 610718 501882 610954
rect 501326 610398 501562 610634
rect 501646 610398 501882 610634
rect 501326 574718 501562 574954
rect 501646 574718 501882 574954
rect 501326 574398 501562 574634
rect 501646 574398 501882 574634
rect 501326 538718 501562 538954
rect 501646 538718 501882 538954
rect 501326 538398 501562 538634
rect 501646 538398 501882 538634
rect 501326 502718 501562 502954
rect 501646 502718 501882 502954
rect 501326 502398 501562 502634
rect 501646 502398 501882 502634
rect 501326 466718 501562 466954
rect 501646 466718 501882 466954
rect 501326 466398 501562 466634
rect 501646 466398 501882 466634
rect 501326 430718 501562 430954
rect 501646 430718 501882 430954
rect 501326 430398 501562 430634
rect 501646 430398 501882 430634
rect 501326 394718 501562 394954
rect 501646 394718 501882 394954
rect 501326 394398 501562 394634
rect 501646 394398 501882 394634
rect 501326 358718 501562 358954
rect 501646 358718 501882 358954
rect 501326 358398 501562 358634
rect 501646 358398 501882 358634
rect 501326 322718 501562 322954
rect 501646 322718 501882 322954
rect 501326 322398 501562 322634
rect 501646 322398 501882 322634
rect 501326 286718 501562 286954
rect 501646 286718 501882 286954
rect 501326 286398 501562 286634
rect 501646 286398 501882 286634
rect 501326 250718 501562 250954
rect 501646 250718 501882 250954
rect 501326 250398 501562 250634
rect 501646 250398 501882 250634
rect 501326 214718 501562 214954
rect 501646 214718 501882 214954
rect 501326 214398 501562 214634
rect 501646 214398 501882 214634
rect 501326 178718 501562 178954
rect 501646 178718 501882 178954
rect 501326 178398 501562 178634
rect 501646 178398 501882 178634
rect 501326 142718 501562 142954
rect 501646 142718 501882 142954
rect 501326 142398 501562 142634
rect 501646 142398 501882 142634
rect 501326 106718 501562 106954
rect 501646 106718 501882 106954
rect 501326 106398 501562 106634
rect 501646 106398 501882 106634
rect 501326 70718 501562 70954
rect 501646 70718 501882 70954
rect 501326 70398 501562 70634
rect 501646 70398 501882 70634
rect 501326 34718 501562 34954
rect 501646 34718 501882 34954
rect 501326 34398 501562 34634
rect 501646 34398 501882 34634
rect 501326 -7302 501562 -7066
rect 501646 -7302 501882 -7066
rect 501326 -7622 501562 -7386
rect 501646 -7622 501882 -7386
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 505826 651218 506062 651454
rect 506146 651218 506382 651454
rect 505826 650898 506062 651134
rect 506146 650898 506382 651134
rect 505826 615218 506062 615454
rect 506146 615218 506382 615454
rect 505826 614898 506062 615134
rect 506146 614898 506382 615134
rect 505826 579218 506062 579454
rect 506146 579218 506382 579454
rect 505826 578898 506062 579134
rect 506146 578898 506382 579134
rect 505826 543218 506062 543454
rect 506146 543218 506382 543454
rect 505826 542898 506062 543134
rect 506146 542898 506382 543134
rect 505826 507218 506062 507454
rect 506146 507218 506382 507454
rect 505826 506898 506062 507134
rect 506146 506898 506382 507134
rect 505826 471218 506062 471454
rect 506146 471218 506382 471454
rect 505826 470898 506062 471134
rect 506146 470898 506382 471134
rect 505826 435218 506062 435454
rect 506146 435218 506382 435454
rect 505826 434898 506062 435134
rect 506146 434898 506382 435134
rect 505826 399218 506062 399454
rect 506146 399218 506382 399454
rect 505826 398898 506062 399134
rect 506146 398898 506382 399134
rect 505826 363218 506062 363454
rect 506146 363218 506382 363454
rect 505826 362898 506062 363134
rect 506146 362898 506382 363134
rect 505826 327218 506062 327454
rect 506146 327218 506382 327454
rect 505826 326898 506062 327134
rect 506146 326898 506382 327134
rect 505826 291218 506062 291454
rect 506146 291218 506382 291454
rect 505826 290898 506062 291134
rect 506146 290898 506382 291134
rect 505826 255218 506062 255454
rect 506146 255218 506382 255454
rect 505826 254898 506062 255134
rect 506146 254898 506382 255134
rect 505826 219218 506062 219454
rect 506146 219218 506382 219454
rect 505826 218898 506062 219134
rect 506146 218898 506382 219134
rect 505826 183218 506062 183454
rect 506146 183218 506382 183454
rect 505826 182898 506062 183134
rect 506146 182898 506382 183134
rect 505826 147218 506062 147454
rect 506146 147218 506382 147454
rect 505826 146898 506062 147134
rect 506146 146898 506382 147134
rect 505826 111218 506062 111454
rect 506146 111218 506382 111454
rect 505826 110898 506062 111134
rect 506146 110898 506382 111134
rect 505826 75218 506062 75454
rect 506146 75218 506382 75454
rect 505826 74898 506062 75134
rect 506146 74898 506382 75134
rect 505826 39218 506062 39454
rect 506146 39218 506382 39454
rect 505826 38898 506062 39134
rect 506146 38898 506382 39134
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 510326 705562 510562 705798
rect 510646 705562 510882 705798
rect 510326 705242 510562 705478
rect 510646 705242 510882 705478
rect 510326 691718 510562 691954
rect 510646 691718 510882 691954
rect 510326 691398 510562 691634
rect 510646 691398 510882 691634
rect 510326 655718 510562 655954
rect 510646 655718 510882 655954
rect 510326 655398 510562 655634
rect 510646 655398 510882 655634
rect 510326 619718 510562 619954
rect 510646 619718 510882 619954
rect 510326 619398 510562 619634
rect 510646 619398 510882 619634
rect 510326 583718 510562 583954
rect 510646 583718 510882 583954
rect 510326 583398 510562 583634
rect 510646 583398 510882 583634
rect 510326 547718 510562 547954
rect 510646 547718 510882 547954
rect 510326 547398 510562 547634
rect 510646 547398 510882 547634
rect 510326 511718 510562 511954
rect 510646 511718 510882 511954
rect 510326 511398 510562 511634
rect 510646 511398 510882 511634
rect 510326 475718 510562 475954
rect 510646 475718 510882 475954
rect 510326 475398 510562 475634
rect 510646 475398 510882 475634
rect 510326 439718 510562 439954
rect 510646 439718 510882 439954
rect 510326 439398 510562 439634
rect 510646 439398 510882 439634
rect 510326 403718 510562 403954
rect 510646 403718 510882 403954
rect 510326 403398 510562 403634
rect 510646 403398 510882 403634
rect 510326 367718 510562 367954
rect 510646 367718 510882 367954
rect 510326 367398 510562 367634
rect 510646 367398 510882 367634
rect 510326 331718 510562 331954
rect 510646 331718 510882 331954
rect 510326 331398 510562 331634
rect 510646 331398 510882 331634
rect 510326 295718 510562 295954
rect 510646 295718 510882 295954
rect 510326 295398 510562 295634
rect 510646 295398 510882 295634
rect 510326 259718 510562 259954
rect 510646 259718 510882 259954
rect 510326 259398 510562 259634
rect 510646 259398 510882 259634
rect 510326 223718 510562 223954
rect 510646 223718 510882 223954
rect 510326 223398 510562 223634
rect 510646 223398 510882 223634
rect 510326 187718 510562 187954
rect 510646 187718 510882 187954
rect 510326 187398 510562 187634
rect 510646 187398 510882 187634
rect 510326 151718 510562 151954
rect 510646 151718 510882 151954
rect 510326 151398 510562 151634
rect 510646 151398 510882 151634
rect 510326 115718 510562 115954
rect 510646 115718 510882 115954
rect 510326 115398 510562 115634
rect 510646 115398 510882 115634
rect 510326 79718 510562 79954
rect 510646 79718 510882 79954
rect 510326 79398 510562 79634
rect 510646 79398 510882 79634
rect 510326 43718 510562 43954
rect 510646 43718 510882 43954
rect 510326 43398 510562 43634
rect 510646 43398 510882 43634
rect 510326 7718 510562 7954
rect 510646 7718 510882 7954
rect 510326 7398 510562 7634
rect 510646 7398 510882 7634
rect 510326 -1542 510562 -1306
rect 510646 -1542 510882 -1306
rect 510326 -1862 510562 -1626
rect 510646 -1862 510882 -1626
rect 514826 706522 515062 706758
rect 515146 706522 515382 706758
rect 514826 706202 515062 706438
rect 515146 706202 515382 706438
rect 514826 696218 515062 696454
rect 515146 696218 515382 696454
rect 514826 695898 515062 696134
rect 515146 695898 515382 696134
rect 514826 660218 515062 660454
rect 515146 660218 515382 660454
rect 514826 659898 515062 660134
rect 515146 659898 515382 660134
rect 514826 624218 515062 624454
rect 515146 624218 515382 624454
rect 514826 623898 515062 624134
rect 515146 623898 515382 624134
rect 514826 588218 515062 588454
rect 515146 588218 515382 588454
rect 514826 587898 515062 588134
rect 515146 587898 515382 588134
rect 514826 552218 515062 552454
rect 515146 552218 515382 552454
rect 514826 551898 515062 552134
rect 515146 551898 515382 552134
rect 514826 516218 515062 516454
rect 515146 516218 515382 516454
rect 514826 515898 515062 516134
rect 515146 515898 515382 516134
rect 514826 480218 515062 480454
rect 515146 480218 515382 480454
rect 514826 479898 515062 480134
rect 515146 479898 515382 480134
rect 514826 444218 515062 444454
rect 515146 444218 515382 444454
rect 514826 443898 515062 444134
rect 515146 443898 515382 444134
rect 514826 408218 515062 408454
rect 515146 408218 515382 408454
rect 514826 407898 515062 408134
rect 515146 407898 515382 408134
rect 514826 372218 515062 372454
rect 515146 372218 515382 372454
rect 514826 371898 515062 372134
rect 515146 371898 515382 372134
rect 514826 336218 515062 336454
rect 515146 336218 515382 336454
rect 514826 335898 515062 336134
rect 515146 335898 515382 336134
rect 514826 300218 515062 300454
rect 515146 300218 515382 300454
rect 514826 299898 515062 300134
rect 515146 299898 515382 300134
rect 514826 264218 515062 264454
rect 515146 264218 515382 264454
rect 514826 263898 515062 264134
rect 515146 263898 515382 264134
rect 514826 228218 515062 228454
rect 515146 228218 515382 228454
rect 514826 227898 515062 228134
rect 515146 227898 515382 228134
rect 514826 192218 515062 192454
rect 515146 192218 515382 192454
rect 514826 191898 515062 192134
rect 515146 191898 515382 192134
rect 514826 156218 515062 156454
rect 515146 156218 515382 156454
rect 514826 155898 515062 156134
rect 515146 155898 515382 156134
rect 514826 120218 515062 120454
rect 515146 120218 515382 120454
rect 514826 119898 515062 120134
rect 515146 119898 515382 120134
rect 514826 84218 515062 84454
rect 515146 84218 515382 84454
rect 514826 83898 515062 84134
rect 515146 83898 515382 84134
rect 514826 48218 515062 48454
rect 515146 48218 515382 48454
rect 514826 47898 515062 48134
rect 515146 47898 515382 48134
rect 514826 12218 515062 12454
rect 515146 12218 515382 12454
rect 514826 11898 515062 12134
rect 515146 11898 515382 12134
rect 514826 -2502 515062 -2266
rect 515146 -2502 515382 -2266
rect 514826 -2822 515062 -2586
rect 515146 -2822 515382 -2586
rect 519326 707482 519562 707718
rect 519646 707482 519882 707718
rect 519326 707162 519562 707398
rect 519646 707162 519882 707398
rect 519326 700718 519562 700954
rect 519646 700718 519882 700954
rect 519326 700398 519562 700634
rect 519646 700398 519882 700634
rect 519326 664718 519562 664954
rect 519646 664718 519882 664954
rect 519326 664398 519562 664634
rect 519646 664398 519882 664634
rect 519326 628718 519562 628954
rect 519646 628718 519882 628954
rect 519326 628398 519562 628634
rect 519646 628398 519882 628634
rect 519326 592718 519562 592954
rect 519646 592718 519882 592954
rect 519326 592398 519562 592634
rect 519646 592398 519882 592634
rect 519326 556718 519562 556954
rect 519646 556718 519882 556954
rect 519326 556398 519562 556634
rect 519646 556398 519882 556634
rect 519326 520718 519562 520954
rect 519646 520718 519882 520954
rect 519326 520398 519562 520634
rect 519646 520398 519882 520634
rect 519326 484718 519562 484954
rect 519646 484718 519882 484954
rect 519326 484398 519562 484634
rect 519646 484398 519882 484634
rect 519326 448718 519562 448954
rect 519646 448718 519882 448954
rect 519326 448398 519562 448634
rect 519646 448398 519882 448634
rect 519326 412718 519562 412954
rect 519646 412718 519882 412954
rect 519326 412398 519562 412634
rect 519646 412398 519882 412634
rect 519326 376718 519562 376954
rect 519646 376718 519882 376954
rect 519326 376398 519562 376634
rect 519646 376398 519882 376634
rect 519326 340718 519562 340954
rect 519646 340718 519882 340954
rect 519326 340398 519562 340634
rect 519646 340398 519882 340634
rect 519326 304718 519562 304954
rect 519646 304718 519882 304954
rect 519326 304398 519562 304634
rect 519646 304398 519882 304634
rect 519326 268718 519562 268954
rect 519646 268718 519882 268954
rect 519326 268398 519562 268634
rect 519646 268398 519882 268634
rect 519326 232718 519562 232954
rect 519646 232718 519882 232954
rect 519326 232398 519562 232634
rect 519646 232398 519882 232634
rect 519326 196718 519562 196954
rect 519646 196718 519882 196954
rect 519326 196398 519562 196634
rect 519646 196398 519882 196634
rect 519326 160718 519562 160954
rect 519646 160718 519882 160954
rect 519326 160398 519562 160634
rect 519646 160398 519882 160634
rect 519326 124718 519562 124954
rect 519646 124718 519882 124954
rect 519326 124398 519562 124634
rect 519646 124398 519882 124634
rect 519326 88718 519562 88954
rect 519646 88718 519882 88954
rect 519326 88398 519562 88634
rect 519646 88398 519882 88634
rect 519326 52718 519562 52954
rect 519646 52718 519882 52954
rect 519326 52398 519562 52634
rect 519646 52398 519882 52634
rect 519326 16718 519562 16954
rect 519646 16718 519882 16954
rect 519326 16398 519562 16634
rect 519646 16398 519882 16634
rect 519326 -3462 519562 -3226
rect 519646 -3462 519882 -3226
rect 519326 -3782 519562 -3546
rect 519646 -3782 519882 -3546
rect 523826 708442 524062 708678
rect 524146 708442 524382 708678
rect 523826 708122 524062 708358
rect 524146 708122 524382 708358
rect 523826 669218 524062 669454
rect 524146 669218 524382 669454
rect 523826 668898 524062 669134
rect 524146 668898 524382 669134
rect 523826 633218 524062 633454
rect 524146 633218 524382 633454
rect 523826 632898 524062 633134
rect 524146 632898 524382 633134
rect 523826 597218 524062 597454
rect 524146 597218 524382 597454
rect 523826 596898 524062 597134
rect 524146 596898 524382 597134
rect 523826 561218 524062 561454
rect 524146 561218 524382 561454
rect 523826 560898 524062 561134
rect 524146 560898 524382 561134
rect 523826 525218 524062 525454
rect 524146 525218 524382 525454
rect 523826 524898 524062 525134
rect 524146 524898 524382 525134
rect 523826 489218 524062 489454
rect 524146 489218 524382 489454
rect 523826 488898 524062 489134
rect 524146 488898 524382 489134
rect 523826 453218 524062 453454
rect 524146 453218 524382 453454
rect 523826 452898 524062 453134
rect 524146 452898 524382 453134
rect 523826 417218 524062 417454
rect 524146 417218 524382 417454
rect 523826 416898 524062 417134
rect 524146 416898 524382 417134
rect 523826 381218 524062 381454
rect 524146 381218 524382 381454
rect 523826 380898 524062 381134
rect 524146 380898 524382 381134
rect 523826 345218 524062 345454
rect 524146 345218 524382 345454
rect 523826 344898 524062 345134
rect 524146 344898 524382 345134
rect 523826 309218 524062 309454
rect 524146 309218 524382 309454
rect 523826 308898 524062 309134
rect 524146 308898 524382 309134
rect 523826 273218 524062 273454
rect 524146 273218 524382 273454
rect 523826 272898 524062 273134
rect 524146 272898 524382 273134
rect 523826 237218 524062 237454
rect 524146 237218 524382 237454
rect 523826 236898 524062 237134
rect 524146 236898 524382 237134
rect 523826 201218 524062 201454
rect 524146 201218 524382 201454
rect 523826 200898 524062 201134
rect 524146 200898 524382 201134
rect 523826 165218 524062 165454
rect 524146 165218 524382 165454
rect 523826 164898 524062 165134
rect 524146 164898 524382 165134
rect 523826 129218 524062 129454
rect 524146 129218 524382 129454
rect 523826 128898 524062 129134
rect 524146 128898 524382 129134
rect 523826 93218 524062 93454
rect 524146 93218 524382 93454
rect 523826 92898 524062 93134
rect 524146 92898 524382 93134
rect 523826 57218 524062 57454
rect 524146 57218 524382 57454
rect 523826 56898 524062 57134
rect 524146 56898 524382 57134
rect 523826 21218 524062 21454
rect 524146 21218 524382 21454
rect 523826 20898 524062 21134
rect 524146 20898 524382 21134
rect 523826 -4422 524062 -4186
rect 524146 -4422 524382 -4186
rect 523826 -4742 524062 -4506
rect 524146 -4742 524382 -4506
rect 528326 709402 528562 709638
rect 528646 709402 528882 709638
rect 528326 709082 528562 709318
rect 528646 709082 528882 709318
rect 528326 673718 528562 673954
rect 528646 673718 528882 673954
rect 528326 673398 528562 673634
rect 528646 673398 528882 673634
rect 528326 637718 528562 637954
rect 528646 637718 528882 637954
rect 528326 637398 528562 637634
rect 528646 637398 528882 637634
rect 528326 601718 528562 601954
rect 528646 601718 528882 601954
rect 528326 601398 528562 601634
rect 528646 601398 528882 601634
rect 528326 565718 528562 565954
rect 528646 565718 528882 565954
rect 528326 565398 528562 565634
rect 528646 565398 528882 565634
rect 528326 529718 528562 529954
rect 528646 529718 528882 529954
rect 528326 529398 528562 529634
rect 528646 529398 528882 529634
rect 528326 493718 528562 493954
rect 528646 493718 528882 493954
rect 528326 493398 528562 493634
rect 528646 493398 528882 493634
rect 528326 457718 528562 457954
rect 528646 457718 528882 457954
rect 528326 457398 528562 457634
rect 528646 457398 528882 457634
rect 528326 421718 528562 421954
rect 528646 421718 528882 421954
rect 528326 421398 528562 421634
rect 528646 421398 528882 421634
rect 528326 385718 528562 385954
rect 528646 385718 528882 385954
rect 528326 385398 528562 385634
rect 528646 385398 528882 385634
rect 528326 349718 528562 349954
rect 528646 349718 528882 349954
rect 528326 349398 528562 349634
rect 528646 349398 528882 349634
rect 528326 313718 528562 313954
rect 528646 313718 528882 313954
rect 528326 313398 528562 313634
rect 528646 313398 528882 313634
rect 528326 277718 528562 277954
rect 528646 277718 528882 277954
rect 528326 277398 528562 277634
rect 528646 277398 528882 277634
rect 528326 241718 528562 241954
rect 528646 241718 528882 241954
rect 528326 241398 528562 241634
rect 528646 241398 528882 241634
rect 528326 205718 528562 205954
rect 528646 205718 528882 205954
rect 528326 205398 528562 205634
rect 528646 205398 528882 205634
rect 528326 169718 528562 169954
rect 528646 169718 528882 169954
rect 528326 169398 528562 169634
rect 528646 169398 528882 169634
rect 528326 133718 528562 133954
rect 528646 133718 528882 133954
rect 528326 133398 528562 133634
rect 528646 133398 528882 133634
rect 528326 97718 528562 97954
rect 528646 97718 528882 97954
rect 528326 97398 528562 97634
rect 528646 97398 528882 97634
rect 528326 61718 528562 61954
rect 528646 61718 528882 61954
rect 528326 61398 528562 61634
rect 528646 61398 528882 61634
rect 528326 25718 528562 25954
rect 528646 25718 528882 25954
rect 528326 25398 528562 25634
rect 528646 25398 528882 25634
rect 528326 -5382 528562 -5146
rect 528646 -5382 528882 -5146
rect 528326 -5702 528562 -5466
rect 528646 -5702 528882 -5466
rect 532826 710362 533062 710598
rect 533146 710362 533382 710598
rect 532826 710042 533062 710278
rect 533146 710042 533382 710278
rect 532826 678218 533062 678454
rect 533146 678218 533382 678454
rect 532826 677898 533062 678134
rect 533146 677898 533382 678134
rect 532826 642218 533062 642454
rect 533146 642218 533382 642454
rect 532826 641898 533062 642134
rect 533146 641898 533382 642134
rect 532826 606218 533062 606454
rect 533146 606218 533382 606454
rect 532826 605898 533062 606134
rect 533146 605898 533382 606134
rect 532826 570218 533062 570454
rect 533146 570218 533382 570454
rect 532826 569898 533062 570134
rect 533146 569898 533382 570134
rect 532826 534218 533062 534454
rect 533146 534218 533382 534454
rect 532826 533898 533062 534134
rect 533146 533898 533382 534134
rect 532826 498218 533062 498454
rect 533146 498218 533382 498454
rect 532826 497898 533062 498134
rect 533146 497898 533382 498134
rect 532826 462218 533062 462454
rect 533146 462218 533382 462454
rect 532826 461898 533062 462134
rect 533146 461898 533382 462134
rect 532826 426218 533062 426454
rect 533146 426218 533382 426454
rect 532826 425898 533062 426134
rect 533146 425898 533382 426134
rect 532826 390218 533062 390454
rect 533146 390218 533382 390454
rect 532826 389898 533062 390134
rect 533146 389898 533382 390134
rect 532826 354218 533062 354454
rect 533146 354218 533382 354454
rect 532826 353898 533062 354134
rect 533146 353898 533382 354134
rect 532826 318218 533062 318454
rect 533146 318218 533382 318454
rect 532826 317898 533062 318134
rect 533146 317898 533382 318134
rect 532826 282218 533062 282454
rect 533146 282218 533382 282454
rect 532826 281898 533062 282134
rect 533146 281898 533382 282134
rect 532826 246218 533062 246454
rect 533146 246218 533382 246454
rect 532826 245898 533062 246134
rect 533146 245898 533382 246134
rect 532826 210218 533062 210454
rect 533146 210218 533382 210454
rect 532826 209898 533062 210134
rect 533146 209898 533382 210134
rect 532826 174218 533062 174454
rect 533146 174218 533382 174454
rect 532826 173898 533062 174134
rect 533146 173898 533382 174134
rect 532826 138218 533062 138454
rect 533146 138218 533382 138454
rect 532826 137898 533062 138134
rect 533146 137898 533382 138134
rect 532826 102218 533062 102454
rect 533146 102218 533382 102454
rect 532826 101898 533062 102134
rect 533146 101898 533382 102134
rect 532826 66218 533062 66454
rect 533146 66218 533382 66454
rect 532826 65898 533062 66134
rect 533146 65898 533382 66134
rect 532826 30218 533062 30454
rect 533146 30218 533382 30454
rect 532826 29898 533062 30134
rect 533146 29898 533382 30134
rect 532826 -6342 533062 -6106
rect 533146 -6342 533382 -6106
rect 532826 -6662 533062 -6426
rect 533146 -6662 533382 -6426
rect 537326 711322 537562 711558
rect 537646 711322 537882 711558
rect 537326 711002 537562 711238
rect 537646 711002 537882 711238
rect 537326 682718 537562 682954
rect 537646 682718 537882 682954
rect 537326 682398 537562 682634
rect 537646 682398 537882 682634
rect 537326 646718 537562 646954
rect 537646 646718 537882 646954
rect 537326 646398 537562 646634
rect 537646 646398 537882 646634
rect 537326 610718 537562 610954
rect 537646 610718 537882 610954
rect 537326 610398 537562 610634
rect 537646 610398 537882 610634
rect 537326 574718 537562 574954
rect 537646 574718 537882 574954
rect 537326 574398 537562 574634
rect 537646 574398 537882 574634
rect 537326 538718 537562 538954
rect 537646 538718 537882 538954
rect 537326 538398 537562 538634
rect 537646 538398 537882 538634
rect 537326 502718 537562 502954
rect 537646 502718 537882 502954
rect 537326 502398 537562 502634
rect 537646 502398 537882 502634
rect 537326 466718 537562 466954
rect 537646 466718 537882 466954
rect 537326 466398 537562 466634
rect 537646 466398 537882 466634
rect 537326 430718 537562 430954
rect 537646 430718 537882 430954
rect 537326 430398 537562 430634
rect 537646 430398 537882 430634
rect 537326 394718 537562 394954
rect 537646 394718 537882 394954
rect 537326 394398 537562 394634
rect 537646 394398 537882 394634
rect 537326 358718 537562 358954
rect 537646 358718 537882 358954
rect 537326 358398 537562 358634
rect 537646 358398 537882 358634
rect 537326 322718 537562 322954
rect 537646 322718 537882 322954
rect 537326 322398 537562 322634
rect 537646 322398 537882 322634
rect 537326 286718 537562 286954
rect 537646 286718 537882 286954
rect 537326 286398 537562 286634
rect 537646 286398 537882 286634
rect 537326 250718 537562 250954
rect 537646 250718 537882 250954
rect 537326 250398 537562 250634
rect 537646 250398 537882 250634
rect 537326 214718 537562 214954
rect 537646 214718 537882 214954
rect 537326 214398 537562 214634
rect 537646 214398 537882 214634
rect 537326 178718 537562 178954
rect 537646 178718 537882 178954
rect 537326 178398 537562 178634
rect 537646 178398 537882 178634
rect 537326 142718 537562 142954
rect 537646 142718 537882 142954
rect 537326 142398 537562 142634
rect 537646 142398 537882 142634
rect 537326 106718 537562 106954
rect 537646 106718 537882 106954
rect 537326 106398 537562 106634
rect 537646 106398 537882 106634
rect 537326 70718 537562 70954
rect 537646 70718 537882 70954
rect 537326 70398 537562 70634
rect 537646 70398 537882 70634
rect 537326 34718 537562 34954
rect 537646 34718 537882 34954
rect 537326 34398 537562 34634
rect 537646 34398 537882 34634
rect 537326 -7302 537562 -7066
rect 537646 -7302 537882 -7066
rect 537326 -7622 537562 -7386
rect 537646 -7622 537882 -7386
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 541826 651218 542062 651454
rect 542146 651218 542382 651454
rect 541826 650898 542062 651134
rect 542146 650898 542382 651134
rect 541826 615218 542062 615454
rect 542146 615218 542382 615454
rect 541826 614898 542062 615134
rect 542146 614898 542382 615134
rect 541826 579218 542062 579454
rect 542146 579218 542382 579454
rect 541826 578898 542062 579134
rect 542146 578898 542382 579134
rect 541826 543218 542062 543454
rect 542146 543218 542382 543454
rect 541826 542898 542062 543134
rect 542146 542898 542382 543134
rect 541826 507218 542062 507454
rect 542146 507218 542382 507454
rect 541826 506898 542062 507134
rect 542146 506898 542382 507134
rect 541826 471218 542062 471454
rect 542146 471218 542382 471454
rect 541826 470898 542062 471134
rect 542146 470898 542382 471134
rect 541826 435218 542062 435454
rect 542146 435218 542382 435454
rect 541826 434898 542062 435134
rect 542146 434898 542382 435134
rect 541826 399218 542062 399454
rect 542146 399218 542382 399454
rect 541826 398898 542062 399134
rect 542146 398898 542382 399134
rect 541826 363218 542062 363454
rect 542146 363218 542382 363454
rect 541826 362898 542062 363134
rect 542146 362898 542382 363134
rect 541826 327218 542062 327454
rect 542146 327218 542382 327454
rect 541826 326898 542062 327134
rect 542146 326898 542382 327134
rect 541826 291218 542062 291454
rect 542146 291218 542382 291454
rect 541826 290898 542062 291134
rect 542146 290898 542382 291134
rect 541826 255218 542062 255454
rect 542146 255218 542382 255454
rect 541826 254898 542062 255134
rect 542146 254898 542382 255134
rect 541826 219218 542062 219454
rect 542146 219218 542382 219454
rect 541826 218898 542062 219134
rect 542146 218898 542382 219134
rect 541826 183218 542062 183454
rect 542146 183218 542382 183454
rect 541826 182898 542062 183134
rect 542146 182898 542382 183134
rect 541826 147218 542062 147454
rect 542146 147218 542382 147454
rect 541826 146898 542062 147134
rect 542146 146898 542382 147134
rect 541826 111218 542062 111454
rect 542146 111218 542382 111454
rect 541826 110898 542062 111134
rect 542146 110898 542382 111134
rect 541826 75218 542062 75454
rect 542146 75218 542382 75454
rect 541826 74898 542062 75134
rect 542146 74898 542382 75134
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 546326 705562 546562 705798
rect 546646 705562 546882 705798
rect 546326 705242 546562 705478
rect 546646 705242 546882 705478
rect 546326 691718 546562 691954
rect 546646 691718 546882 691954
rect 546326 691398 546562 691634
rect 546646 691398 546882 691634
rect 546326 655718 546562 655954
rect 546646 655718 546882 655954
rect 546326 655398 546562 655634
rect 546646 655398 546882 655634
rect 546326 619718 546562 619954
rect 546646 619718 546882 619954
rect 546326 619398 546562 619634
rect 546646 619398 546882 619634
rect 546326 583718 546562 583954
rect 546646 583718 546882 583954
rect 546326 583398 546562 583634
rect 546646 583398 546882 583634
rect 546326 547718 546562 547954
rect 546646 547718 546882 547954
rect 546326 547398 546562 547634
rect 546646 547398 546882 547634
rect 546326 511718 546562 511954
rect 546646 511718 546882 511954
rect 546326 511398 546562 511634
rect 546646 511398 546882 511634
rect 546326 475718 546562 475954
rect 546646 475718 546882 475954
rect 546326 475398 546562 475634
rect 546646 475398 546882 475634
rect 546326 439718 546562 439954
rect 546646 439718 546882 439954
rect 546326 439398 546562 439634
rect 546646 439398 546882 439634
rect 546326 403718 546562 403954
rect 546646 403718 546882 403954
rect 546326 403398 546562 403634
rect 546646 403398 546882 403634
rect 546326 367718 546562 367954
rect 546646 367718 546882 367954
rect 546326 367398 546562 367634
rect 546646 367398 546882 367634
rect 546326 331718 546562 331954
rect 546646 331718 546882 331954
rect 546326 331398 546562 331634
rect 546646 331398 546882 331634
rect 546326 295718 546562 295954
rect 546646 295718 546882 295954
rect 546326 295398 546562 295634
rect 546646 295398 546882 295634
rect 546326 259718 546562 259954
rect 546646 259718 546882 259954
rect 546326 259398 546562 259634
rect 546646 259398 546882 259634
rect 546326 223718 546562 223954
rect 546646 223718 546882 223954
rect 546326 223398 546562 223634
rect 546646 223398 546882 223634
rect 546326 187718 546562 187954
rect 546646 187718 546882 187954
rect 546326 187398 546562 187634
rect 546646 187398 546882 187634
rect 546326 151718 546562 151954
rect 546646 151718 546882 151954
rect 546326 151398 546562 151634
rect 546646 151398 546882 151634
rect 546326 115718 546562 115954
rect 546646 115718 546882 115954
rect 546326 115398 546562 115634
rect 546646 115398 546882 115634
rect 546326 79718 546562 79954
rect 546646 79718 546882 79954
rect 546326 79398 546562 79634
rect 546646 79398 546882 79634
rect 546326 43718 546562 43954
rect 546646 43718 546882 43954
rect 546326 43398 546562 43634
rect 546646 43398 546882 43634
rect 546326 7718 546562 7954
rect 546646 7718 546882 7954
rect 546326 7398 546562 7634
rect 546646 7398 546882 7634
rect 546326 -1542 546562 -1306
rect 546646 -1542 546882 -1306
rect 546326 -1862 546562 -1626
rect 546646 -1862 546882 -1626
rect 550826 706522 551062 706758
rect 551146 706522 551382 706758
rect 550826 706202 551062 706438
rect 551146 706202 551382 706438
rect 550826 696218 551062 696454
rect 551146 696218 551382 696454
rect 550826 695898 551062 696134
rect 551146 695898 551382 696134
rect 550826 660218 551062 660454
rect 551146 660218 551382 660454
rect 550826 659898 551062 660134
rect 551146 659898 551382 660134
rect 550826 624218 551062 624454
rect 551146 624218 551382 624454
rect 550826 623898 551062 624134
rect 551146 623898 551382 624134
rect 550826 588218 551062 588454
rect 551146 588218 551382 588454
rect 550826 587898 551062 588134
rect 551146 587898 551382 588134
rect 550826 552218 551062 552454
rect 551146 552218 551382 552454
rect 550826 551898 551062 552134
rect 551146 551898 551382 552134
rect 550826 516218 551062 516454
rect 551146 516218 551382 516454
rect 550826 515898 551062 516134
rect 551146 515898 551382 516134
rect 550826 480218 551062 480454
rect 551146 480218 551382 480454
rect 550826 479898 551062 480134
rect 551146 479898 551382 480134
rect 550826 444218 551062 444454
rect 551146 444218 551382 444454
rect 550826 443898 551062 444134
rect 551146 443898 551382 444134
rect 550826 408218 551062 408454
rect 551146 408218 551382 408454
rect 550826 407898 551062 408134
rect 551146 407898 551382 408134
rect 550826 372218 551062 372454
rect 551146 372218 551382 372454
rect 550826 371898 551062 372134
rect 551146 371898 551382 372134
rect 550826 336218 551062 336454
rect 551146 336218 551382 336454
rect 550826 335898 551062 336134
rect 551146 335898 551382 336134
rect 550826 300218 551062 300454
rect 551146 300218 551382 300454
rect 550826 299898 551062 300134
rect 551146 299898 551382 300134
rect 550826 264218 551062 264454
rect 551146 264218 551382 264454
rect 550826 263898 551062 264134
rect 551146 263898 551382 264134
rect 550826 228218 551062 228454
rect 551146 228218 551382 228454
rect 550826 227898 551062 228134
rect 551146 227898 551382 228134
rect 550826 192218 551062 192454
rect 551146 192218 551382 192454
rect 550826 191898 551062 192134
rect 551146 191898 551382 192134
rect 550826 156218 551062 156454
rect 551146 156218 551382 156454
rect 550826 155898 551062 156134
rect 551146 155898 551382 156134
rect 550826 120218 551062 120454
rect 551146 120218 551382 120454
rect 550826 119898 551062 120134
rect 551146 119898 551382 120134
rect 550826 84218 551062 84454
rect 551146 84218 551382 84454
rect 550826 83898 551062 84134
rect 551146 83898 551382 84134
rect 550826 48218 551062 48454
rect 551146 48218 551382 48454
rect 550826 47898 551062 48134
rect 551146 47898 551382 48134
rect 550826 12218 551062 12454
rect 551146 12218 551382 12454
rect 550826 11898 551062 12134
rect 551146 11898 551382 12134
rect 550826 -2502 551062 -2266
rect 551146 -2502 551382 -2266
rect 550826 -2822 551062 -2586
rect 551146 -2822 551382 -2586
rect 555326 707482 555562 707718
rect 555646 707482 555882 707718
rect 555326 707162 555562 707398
rect 555646 707162 555882 707398
rect 555326 700718 555562 700954
rect 555646 700718 555882 700954
rect 555326 700398 555562 700634
rect 555646 700398 555882 700634
rect 555326 664718 555562 664954
rect 555646 664718 555882 664954
rect 555326 664398 555562 664634
rect 555646 664398 555882 664634
rect 555326 628718 555562 628954
rect 555646 628718 555882 628954
rect 555326 628398 555562 628634
rect 555646 628398 555882 628634
rect 555326 592718 555562 592954
rect 555646 592718 555882 592954
rect 555326 592398 555562 592634
rect 555646 592398 555882 592634
rect 555326 556718 555562 556954
rect 555646 556718 555882 556954
rect 555326 556398 555562 556634
rect 555646 556398 555882 556634
rect 555326 520718 555562 520954
rect 555646 520718 555882 520954
rect 555326 520398 555562 520634
rect 555646 520398 555882 520634
rect 555326 484718 555562 484954
rect 555646 484718 555882 484954
rect 555326 484398 555562 484634
rect 555646 484398 555882 484634
rect 555326 448718 555562 448954
rect 555646 448718 555882 448954
rect 555326 448398 555562 448634
rect 555646 448398 555882 448634
rect 555326 412718 555562 412954
rect 555646 412718 555882 412954
rect 555326 412398 555562 412634
rect 555646 412398 555882 412634
rect 555326 376718 555562 376954
rect 555646 376718 555882 376954
rect 555326 376398 555562 376634
rect 555646 376398 555882 376634
rect 555326 340718 555562 340954
rect 555646 340718 555882 340954
rect 555326 340398 555562 340634
rect 555646 340398 555882 340634
rect 555326 304718 555562 304954
rect 555646 304718 555882 304954
rect 555326 304398 555562 304634
rect 555646 304398 555882 304634
rect 555326 268718 555562 268954
rect 555646 268718 555882 268954
rect 555326 268398 555562 268634
rect 555646 268398 555882 268634
rect 555326 232718 555562 232954
rect 555646 232718 555882 232954
rect 555326 232398 555562 232634
rect 555646 232398 555882 232634
rect 555326 196718 555562 196954
rect 555646 196718 555882 196954
rect 555326 196398 555562 196634
rect 555646 196398 555882 196634
rect 555326 160718 555562 160954
rect 555646 160718 555882 160954
rect 555326 160398 555562 160634
rect 555646 160398 555882 160634
rect 555326 124718 555562 124954
rect 555646 124718 555882 124954
rect 555326 124398 555562 124634
rect 555646 124398 555882 124634
rect 555326 88718 555562 88954
rect 555646 88718 555882 88954
rect 555326 88398 555562 88634
rect 555646 88398 555882 88634
rect 555326 52718 555562 52954
rect 555646 52718 555882 52954
rect 555326 52398 555562 52634
rect 555646 52398 555882 52634
rect 555326 16718 555562 16954
rect 555646 16718 555882 16954
rect 555326 16398 555562 16634
rect 555646 16398 555882 16634
rect 555326 -3462 555562 -3226
rect 555646 -3462 555882 -3226
rect 555326 -3782 555562 -3546
rect 555646 -3782 555882 -3546
rect 559826 708442 560062 708678
rect 560146 708442 560382 708678
rect 559826 708122 560062 708358
rect 560146 708122 560382 708358
rect 559826 669218 560062 669454
rect 560146 669218 560382 669454
rect 559826 668898 560062 669134
rect 560146 668898 560382 669134
rect 559826 633218 560062 633454
rect 560146 633218 560382 633454
rect 559826 632898 560062 633134
rect 560146 632898 560382 633134
rect 559826 597218 560062 597454
rect 560146 597218 560382 597454
rect 559826 596898 560062 597134
rect 560146 596898 560382 597134
rect 559826 561218 560062 561454
rect 560146 561218 560382 561454
rect 559826 560898 560062 561134
rect 560146 560898 560382 561134
rect 559826 525218 560062 525454
rect 560146 525218 560382 525454
rect 559826 524898 560062 525134
rect 560146 524898 560382 525134
rect 559826 489218 560062 489454
rect 560146 489218 560382 489454
rect 559826 488898 560062 489134
rect 560146 488898 560382 489134
rect 559826 453218 560062 453454
rect 560146 453218 560382 453454
rect 559826 452898 560062 453134
rect 560146 452898 560382 453134
rect 559826 417218 560062 417454
rect 560146 417218 560382 417454
rect 559826 416898 560062 417134
rect 560146 416898 560382 417134
rect 559826 381218 560062 381454
rect 560146 381218 560382 381454
rect 559826 380898 560062 381134
rect 560146 380898 560382 381134
rect 559826 345218 560062 345454
rect 560146 345218 560382 345454
rect 559826 344898 560062 345134
rect 560146 344898 560382 345134
rect 559826 309218 560062 309454
rect 560146 309218 560382 309454
rect 559826 308898 560062 309134
rect 560146 308898 560382 309134
rect 559826 273218 560062 273454
rect 560146 273218 560382 273454
rect 559826 272898 560062 273134
rect 560146 272898 560382 273134
rect 559826 237218 560062 237454
rect 560146 237218 560382 237454
rect 559826 236898 560062 237134
rect 560146 236898 560382 237134
rect 559826 201218 560062 201454
rect 560146 201218 560382 201454
rect 559826 200898 560062 201134
rect 560146 200898 560382 201134
rect 559826 165218 560062 165454
rect 560146 165218 560382 165454
rect 559826 164898 560062 165134
rect 560146 164898 560382 165134
rect 559826 129218 560062 129454
rect 560146 129218 560382 129454
rect 559826 128898 560062 129134
rect 560146 128898 560382 129134
rect 559826 93218 560062 93454
rect 560146 93218 560382 93454
rect 559826 92898 560062 93134
rect 560146 92898 560382 93134
rect 559826 57218 560062 57454
rect 560146 57218 560382 57454
rect 559826 56898 560062 57134
rect 560146 56898 560382 57134
rect 559826 21218 560062 21454
rect 560146 21218 560382 21454
rect 559826 20898 560062 21134
rect 560146 20898 560382 21134
rect 559826 -4422 560062 -4186
rect 560146 -4422 560382 -4186
rect 559826 -4742 560062 -4506
rect 560146 -4742 560382 -4506
rect 564326 709402 564562 709638
rect 564646 709402 564882 709638
rect 564326 709082 564562 709318
rect 564646 709082 564882 709318
rect 564326 673718 564562 673954
rect 564646 673718 564882 673954
rect 564326 673398 564562 673634
rect 564646 673398 564882 673634
rect 564326 637718 564562 637954
rect 564646 637718 564882 637954
rect 564326 637398 564562 637634
rect 564646 637398 564882 637634
rect 564326 601718 564562 601954
rect 564646 601718 564882 601954
rect 564326 601398 564562 601634
rect 564646 601398 564882 601634
rect 564326 565718 564562 565954
rect 564646 565718 564882 565954
rect 564326 565398 564562 565634
rect 564646 565398 564882 565634
rect 564326 529718 564562 529954
rect 564646 529718 564882 529954
rect 564326 529398 564562 529634
rect 564646 529398 564882 529634
rect 564326 493718 564562 493954
rect 564646 493718 564882 493954
rect 564326 493398 564562 493634
rect 564646 493398 564882 493634
rect 564326 457718 564562 457954
rect 564646 457718 564882 457954
rect 564326 457398 564562 457634
rect 564646 457398 564882 457634
rect 564326 421718 564562 421954
rect 564646 421718 564882 421954
rect 564326 421398 564562 421634
rect 564646 421398 564882 421634
rect 564326 385718 564562 385954
rect 564646 385718 564882 385954
rect 564326 385398 564562 385634
rect 564646 385398 564882 385634
rect 564326 349718 564562 349954
rect 564646 349718 564882 349954
rect 564326 349398 564562 349634
rect 564646 349398 564882 349634
rect 564326 313718 564562 313954
rect 564646 313718 564882 313954
rect 564326 313398 564562 313634
rect 564646 313398 564882 313634
rect 564326 277718 564562 277954
rect 564646 277718 564882 277954
rect 564326 277398 564562 277634
rect 564646 277398 564882 277634
rect 564326 241718 564562 241954
rect 564646 241718 564882 241954
rect 564326 241398 564562 241634
rect 564646 241398 564882 241634
rect 564326 205718 564562 205954
rect 564646 205718 564882 205954
rect 564326 205398 564562 205634
rect 564646 205398 564882 205634
rect 564326 169718 564562 169954
rect 564646 169718 564882 169954
rect 564326 169398 564562 169634
rect 564646 169398 564882 169634
rect 564326 133718 564562 133954
rect 564646 133718 564882 133954
rect 564326 133398 564562 133634
rect 564646 133398 564882 133634
rect 564326 97718 564562 97954
rect 564646 97718 564882 97954
rect 564326 97398 564562 97634
rect 564646 97398 564882 97634
rect 564326 61718 564562 61954
rect 564646 61718 564882 61954
rect 564326 61398 564562 61634
rect 564646 61398 564882 61634
rect 564326 25718 564562 25954
rect 564646 25718 564882 25954
rect 564326 25398 564562 25634
rect 564646 25398 564882 25634
rect 564326 -5382 564562 -5146
rect 564646 -5382 564882 -5146
rect 564326 -5702 564562 -5466
rect 564646 -5702 564882 -5466
rect 568826 710362 569062 710598
rect 569146 710362 569382 710598
rect 568826 710042 569062 710278
rect 569146 710042 569382 710278
rect 568826 678218 569062 678454
rect 569146 678218 569382 678454
rect 568826 677898 569062 678134
rect 569146 677898 569382 678134
rect 568826 642218 569062 642454
rect 569146 642218 569382 642454
rect 568826 641898 569062 642134
rect 569146 641898 569382 642134
rect 568826 606218 569062 606454
rect 569146 606218 569382 606454
rect 568826 605898 569062 606134
rect 569146 605898 569382 606134
rect 568826 570218 569062 570454
rect 569146 570218 569382 570454
rect 568826 569898 569062 570134
rect 569146 569898 569382 570134
rect 568826 534218 569062 534454
rect 569146 534218 569382 534454
rect 568826 533898 569062 534134
rect 569146 533898 569382 534134
rect 568826 498218 569062 498454
rect 569146 498218 569382 498454
rect 568826 497898 569062 498134
rect 569146 497898 569382 498134
rect 568826 462218 569062 462454
rect 569146 462218 569382 462454
rect 568826 461898 569062 462134
rect 569146 461898 569382 462134
rect 568826 426218 569062 426454
rect 569146 426218 569382 426454
rect 568826 425898 569062 426134
rect 569146 425898 569382 426134
rect 568826 390218 569062 390454
rect 569146 390218 569382 390454
rect 568826 389898 569062 390134
rect 569146 389898 569382 390134
rect 568826 354218 569062 354454
rect 569146 354218 569382 354454
rect 568826 353898 569062 354134
rect 569146 353898 569382 354134
rect 568826 318218 569062 318454
rect 569146 318218 569382 318454
rect 568826 317898 569062 318134
rect 569146 317898 569382 318134
rect 568826 282218 569062 282454
rect 569146 282218 569382 282454
rect 568826 281898 569062 282134
rect 569146 281898 569382 282134
rect 568826 246218 569062 246454
rect 569146 246218 569382 246454
rect 568826 245898 569062 246134
rect 569146 245898 569382 246134
rect 568826 210218 569062 210454
rect 569146 210218 569382 210454
rect 568826 209898 569062 210134
rect 569146 209898 569382 210134
rect 568826 174218 569062 174454
rect 569146 174218 569382 174454
rect 568826 173898 569062 174134
rect 569146 173898 569382 174134
rect 568826 138218 569062 138454
rect 569146 138218 569382 138454
rect 568826 137898 569062 138134
rect 569146 137898 569382 138134
rect 568826 102218 569062 102454
rect 569146 102218 569382 102454
rect 568826 101898 569062 102134
rect 569146 101898 569382 102134
rect 568826 66218 569062 66454
rect 569146 66218 569382 66454
rect 568826 65898 569062 66134
rect 569146 65898 569382 66134
rect 568826 30218 569062 30454
rect 569146 30218 569382 30454
rect 568826 29898 569062 30134
rect 569146 29898 569382 30134
rect 568826 -6342 569062 -6106
rect 569146 -6342 569382 -6106
rect 568826 -6662 569062 -6426
rect 569146 -6662 569382 -6426
rect 573326 711322 573562 711558
rect 573646 711322 573882 711558
rect 573326 711002 573562 711238
rect 573646 711002 573882 711238
rect 573326 682718 573562 682954
rect 573646 682718 573882 682954
rect 573326 682398 573562 682634
rect 573646 682398 573882 682634
rect 573326 646718 573562 646954
rect 573646 646718 573882 646954
rect 573326 646398 573562 646634
rect 573646 646398 573882 646634
rect 573326 610718 573562 610954
rect 573646 610718 573882 610954
rect 573326 610398 573562 610634
rect 573646 610398 573882 610634
rect 573326 574718 573562 574954
rect 573646 574718 573882 574954
rect 573326 574398 573562 574634
rect 573646 574398 573882 574634
rect 573326 538718 573562 538954
rect 573646 538718 573882 538954
rect 573326 538398 573562 538634
rect 573646 538398 573882 538634
rect 573326 502718 573562 502954
rect 573646 502718 573882 502954
rect 573326 502398 573562 502634
rect 573646 502398 573882 502634
rect 573326 466718 573562 466954
rect 573646 466718 573882 466954
rect 573326 466398 573562 466634
rect 573646 466398 573882 466634
rect 573326 430718 573562 430954
rect 573646 430718 573882 430954
rect 573326 430398 573562 430634
rect 573646 430398 573882 430634
rect 573326 394718 573562 394954
rect 573646 394718 573882 394954
rect 573326 394398 573562 394634
rect 573646 394398 573882 394634
rect 573326 358718 573562 358954
rect 573646 358718 573882 358954
rect 573326 358398 573562 358634
rect 573646 358398 573882 358634
rect 573326 322718 573562 322954
rect 573646 322718 573882 322954
rect 573326 322398 573562 322634
rect 573646 322398 573882 322634
rect 573326 286718 573562 286954
rect 573646 286718 573882 286954
rect 573326 286398 573562 286634
rect 573646 286398 573882 286634
rect 573326 250718 573562 250954
rect 573646 250718 573882 250954
rect 573326 250398 573562 250634
rect 573646 250398 573882 250634
rect 573326 214718 573562 214954
rect 573646 214718 573882 214954
rect 573326 214398 573562 214634
rect 573646 214398 573882 214634
rect 573326 178718 573562 178954
rect 573646 178718 573882 178954
rect 573326 178398 573562 178634
rect 573646 178398 573882 178634
rect 573326 142718 573562 142954
rect 573646 142718 573882 142954
rect 573326 142398 573562 142634
rect 573646 142398 573882 142634
rect 573326 106718 573562 106954
rect 573646 106718 573882 106954
rect 573326 106398 573562 106634
rect 573646 106398 573882 106634
rect 573326 70718 573562 70954
rect 573646 70718 573882 70954
rect 573326 70398 573562 70634
rect 573646 70398 573882 70634
rect 573326 34718 573562 34954
rect 573646 34718 573882 34954
rect 573326 34398 573562 34634
rect 573646 34398 573882 34634
rect 573326 -7302 573562 -7066
rect 573646 -7302 573882 -7066
rect 573326 -7622 573562 -7386
rect 573646 -7622 573882 -7386
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 582326 705562 582562 705798
rect 582646 705562 582882 705798
rect 582326 705242 582562 705478
rect 582646 705242 582882 705478
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 582326 691718 582562 691954
rect 582646 691718 582882 691954
rect 582326 691398 582562 691634
rect 582646 691398 582882 691634
rect 582326 655718 582562 655954
rect 582646 655718 582882 655954
rect 582326 655398 582562 655634
rect 582646 655398 582882 655634
rect 582326 619718 582562 619954
rect 582646 619718 582882 619954
rect 582326 619398 582562 619634
rect 582646 619398 582882 619634
rect 582326 583718 582562 583954
rect 582646 583718 582882 583954
rect 582326 583398 582562 583634
rect 582646 583398 582882 583634
rect 582326 547718 582562 547954
rect 582646 547718 582882 547954
rect 582326 547398 582562 547634
rect 582646 547398 582882 547634
rect 582326 511718 582562 511954
rect 582646 511718 582882 511954
rect 582326 511398 582562 511634
rect 582646 511398 582882 511634
rect 582326 475718 582562 475954
rect 582646 475718 582882 475954
rect 582326 475398 582562 475634
rect 582646 475398 582882 475634
rect 582326 439718 582562 439954
rect 582646 439718 582882 439954
rect 582326 439398 582562 439634
rect 582646 439398 582882 439634
rect 582326 403718 582562 403954
rect 582646 403718 582882 403954
rect 582326 403398 582562 403634
rect 582646 403398 582882 403634
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 582326 367718 582562 367954
rect 582646 367718 582882 367954
rect 582326 367398 582562 367634
rect 582646 367398 582882 367634
rect 582326 331718 582562 331954
rect 582646 331718 582882 331954
rect 582326 331398 582562 331634
rect 582646 331398 582882 331634
rect 582326 295718 582562 295954
rect 582646 295718 582882 295954
rect 582326 295398 582562 295634
rect 582646 295398 582882 295634
rect 582326 259718 582562 259954
rect 582646 259718 582882 259954
rect 582326 259398 582562 259634
rect 582646 259398 582882 259634
rect 582326 223718 582562 223954
rect 582646 223718 582882 223954
rect 582326 223398 582562 223634
rect 582646 223398 582882 223634
rect 582326 187718 582562 187954
rect 582646 187718 582882 187954
rect 582326 187398 582562 187634
rect 582646 187398 582882 187634
rect 582326 151718 582562 151954
rect 582646 151718 582882 151954
rect 582326 151398 582562 151634
rect 582646 151398 582882 151634
rect 582326 115718 582562 115954
rect 582646 115718 582882 115954
rect 582326 115398 582562 115634
rect 582646 115398 582882 115634
rect 582326 79718 582562 79954
rect 582646 79718 582882 79954
rect 582326 79398 582562 79634
rect 582646 79398 582882 79634
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 582326 43718 582562 43954
rect 582646 43718 582882 43954
rect 582326 43398 582562 43634
rect 582646 43398 582882 43634
rect 582326 7718 582562 7954
rect 582646 7718 582882 7954
rect 582326 7398 582562 7634
rect 582646 7398 582882 7634
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 691718 586538 691954
rect 586622 691718 586858 691954
rect 586302 691398 586538 691634
rect 586622 691398 586858 691634
rect 586302 655718 586538 655954
rect 586622 655718 586858 655954
rect 586302 655398 586538 655634
rect 586622 655398 586858 655634
rect 586302 619718 586538 619954
rect 586622 619718 586858 619954
rect 586302 619398 586538 619634
rect 586622 619398 586858 619634
rect 586302 583718 586538 583954
rect 586622 583718 586858 583954
rect 586302 583398 586538 583634
rect 586622 583398 586858 583634
rect 586302 547718 586538 547954
rect 586622 547718 586858 547954
rect 586302 547398 586538 547634
rect 586622 547398 586858 547634
rect 586302 511718 586538 511954
rect 586622 511718 586858 511954
rect 586302 511398 586538 511634
rect 586622 511398 586858 511634
rect 586302 475718 586538 475954
rect 586622 475718 586858 475954
rect 586302 475398 586538 475634
rect 586622 475398 586858 475634
rect 586302 439718 586538 439954
rect 586622 439718 586858 439954
rect 586302 439398 586538 439634
rect 586622 439398 586858 439634
rect 586302 403718 586538 403954
rect 586622 403718 586858 403954
rect 586302 403398 586538 403634
rect 586622 403398 586858 403634
rect 586302 367718 586538 367954
rect 586622 367718 586858 367954
rect 586302 367398 586538 367634
rect 586622 367398 586858 367634
rect 586302 331718 586538 331954
rect 586622 331718 586858 331954
rect 586302 331398 586538 331634
rect 586622 331398 586858 331634
rect 586302 295718 586538 295954
rect 586622 295718 586858 295954
rect 586302 295398 586538 295634
rect 586622 295398 586858 295634
rect 586302 259718 586538 259954
rect 586622 259718 586858 259954
rect 586302 259398 586538 259634
rect 586622 259398 586858 259634
rect 586302 223718 586538 223954
rect 586622 223718 586858 223954
rect 586302 223398 586538 223634
rect 586622 223398 586858 223634
rect 586302 187718 586538 187954
rect 586622 187718 586858 187954
rect 586302 187398 586538 187634
rect 586622 187398 586858 187634
rect 586302 151718 586538 151954
rect 586622 151718 586858 151954
rect 586302 151398 586538 151634
rect 586622 151398 586858 151634
rect 586302 115718 586538 115954
rect 586622 115718 586858 115954
rect 586302 115398 586538 115634
rect 586622 115398 586858 115634
rect 586302 79718 586538 79954
rect 586622 79718 586858 79954
rect 586302 79398 586538 79634
rect 586622 79398 586858 79634
rect 586302 43718 586538 43954
rect 586622 43718 586858 43954
rect 586302 43398 586538 43634
rect 586622 43398 586858 43634
rect 586302 7718 586538 7954
rect 586622 7718 586858 7954
rect 586302 7398 586538 7634
rect 586622 7398 586858 7634
rect 582326 -1542 582562 -1306
rect 582646 -1542 582882 -1306
rect 582326 -1862 582562 -1626
rect 582646 -1862 582882 -1626
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 696218 587498 696454
rect 587582 696218 587818 696454
rect 587262 695898 587498 696134
rect 587582 695898 587818 696134
rect 587262 660218 587498 660454
rect 587582 660218 587818 660454
rect 587262 659898 587498 660134
rect 587582 659898 587818 660134
rect 587262 624218 587498 624454
rect 587582 624218 587818 624454
rect 587262 623898 587498 624134
rect 587582 623898 587818 624134
rect 587262 588218 587498 588454
rect 587582 588218 587818 588454
rect 587262 587898 587498 588134
rect 587582 587898 587818 588134
rect 587262 552218 587498 552454
rect 587582 552218 587818 552454
rect 587262 551898 587498 552134
rect 587582 551898 587818 552134
rect 587262 516218 587498 516454
rect 587582 516218 587818 516454
rect 587262 515898 587498 516134
rect 587582 515898 587818 516134
rect 587262 480218 587498 480454
rect 587582 480218 587818 480454
rect 587262 479898 587498 480134
rect 587582 479898 587818 480134
rect 587262 444218 587498 444454
rect 587582 444218 587818 444454
rect 587262 443898 587498 444134
rect 587582 443898 587818 444134
rect 587262 408218 587498 408454
rect 587582 408218 587818 408454
rect 587262 407898 587498 408134
rect 587582 407898 587818 408134
rect 587262 372218 587498 372454
rect 587582 372218 587818 372454
rect 587262 371898 587498 372134
rect 587582 371898 587818 372134
rect 587262 336218 587498 336454
rect 587582 336218 587818 336454
rect 587262 335898 587498 336134
rect 587582 335898 587818 336134
rect 587262 300218 587498 300454
rect 587582 300218 587818 300454
rect 587262 299898 587498 300134
rect 587582 299898 587818 300134
rect 587262 264218 587498 264454
rect 587582 264218 587818 264454
rect 587262 263898 587498 264134
rect 587582 263898 587818 264134
rect 587262 228218 587498 228454
rect 587582 228218 587818 228454
rect 587262 227898 587498 228134
rect 587582 227898 587818 228134
rect 587262 192218 587498 192454
rect 587582 192218 587818 192454
rect 587262 191898 587498 192134
rect 587582 191898 587818 192134
rect 587262 156218 587498 156454
rect 587582 156218 587818 156454
rect 587262 155898 587498 156134
rect 587582 155898 587818 156134
rect 587262 120218 587498 120454
rect 587582 120218 587818 120454
rect 587262 119898 587498 120134
rect 587582 119898 587818 120134
rect 587262 84218 587498 84454
rect 587582 84218 587818 84454
rect 587262 83898 587498 84134
rect 587582 83898 587818 84134
rect 587262 48218 587498 48454
rect 587582 48218 587818 48454
rect 587262 47898 587498 48134
rect 587582 47898 587818 48134
rect 587262 12218 587498 12454
rect 587582 12218 587818 12454
rect 587262 11898 587498 12134
rect 587582 11898 587818 12134
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 700718 588458 700954
rect 588542 700718 588778 700954
rect 588222 700398 588458 700634
rect 588542 700398 588778 700634
rect 588222 664718 588458 664954
rect 588542 664718 588778 664954
rect 588222 664398 588458 664634
rect 588542 664398 588778 664634
rect 588222 628718 588458 628954
rect 588542 628718 588778 628954
rect 588222 628398 588458 628634
rect 588542 628398 588778 628634
rect 588222 592718 588458 592954
rect 588542 592718 588778 592954
rect 588222 592398 588458 592634
rect 588542 592398 588778 592634
rect 588222 556718 588458 556954
rect 588542 556718 588778 556954
rect 588222 556398 588458 556634
rect 588542 556398 588778 556634
rect 588222 520718 588458 520954
rect 588542 520718 588778 520954
rect 588222 520398 588458 520634
rect 588542 520398 588778 520634
rect 588222 484718 588458 484954
rect 588542 484718 588778 484954
rect 588222 484398 588458 484634
rect 588542 484398 588778 484634
rect 588222 448718 588458 448954
rect 588542 448718 588778 448954
rect 588222 448398 588458 448634
rect 588542 448398 588778 448634
rect 588222 412718 588458 412954
rect 588542 412718 588778 412954
rect 588222 412398 588458 412634
rect 588542 412398 588778 412634
rect 588222 376718 588458 376954
rect 588542 376718 588778 376954
rect 588222 376398 588458 376634
rect 588542 376398 588778 376634
rect 588222 340718 588458 340954
rect 588542 340718 588778 340954
rect 588222 340398 588458 340634
rect 588542 340398 588778 340634
rect 588222 304718 588458 304954
rect 588542 304718 588778 304954
rect 588222 304398 588458 304634
rect 588542 304398 588778 304634
rect 588222 268718 588458 268954
rect 588542 268718 588778 268954
rect 588222 268398 588458 268634
rect 588542 268398 588778 268634
rect 588222 232718 588458 232954
rect 588542 232718 588778 232954
rect 588222 232398 588458 232634
rect 588542 232398 588778 232634
rect 588222 196718 588458 196954
rect 588542 196718 588778 196954
rect 588222 196398 588458 196634
rect 588542 196398 588778 196634
rect 588222 160718 588458 160954
rect 588542 160718 588778 160954
rect 588222 160398 588458 160634
rect 588542 160398 588778 160634
rect 588222 124718 588458 124954
rect 588542 124718 588778 124954
rect 588222 124398 588458 124634
rect 588542 124398 588778 124634
rect 588222 88718 588458 88954
rect 588542 88718 588778 88954
rect 588222 88398 588458 88634
rect 588542 88398 588778 88634
rect 588222 52718 588458 52954
rect 588542 52718 588778 52954
rect 588222 52398 588458 52634
rect 588542 52398 588778 52634
rect 588222 16718 588458 16954
rect 588542 16718 588778 16954
rect 588222 16398 588458 16634
rect 588542 16398 588778 16634
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 669218 589418 669454
rect 589502 669218 589738 669454
rect 589182 668898 589418 669134
rect 589502 668898 589738 669134
rect 589182 633218 589418 633454
rect 589502 633218 589738 633454
rect 589182 632898 589418 633134
rect 589502 632898 589738 633134
rect 589182 597218 589418 597454
rect 589502 597218 589738 597454
rect 589182 596898 589418 597134
rect 589502 596898 589738 597134
rect 589182 561218 589418 561454
rect 589502 561218 589738 561454
rect 589182 560898 589418 561134
rect 589502 560898 589738 561134
rect 589182 525218 589418 525454
rect 589502 525218 589738 525454
rect 589182 524898 589418 525134
rect 589502 524898 589738 525134
rect 589182 489218 589418 489454
rect 589502 489218 589738 489454
rect 589182 488898 589418 489134
rect 589502 488898 589738 489134
rect 589182 453218 589418 453454
rect 589502 453218 589738 453454
rect 589182 452898 589418 453134
rect 589502 452898 589738 453134
rect 589182 417218 589418 417454
rect 589502 417218 589738 417454
rect 589182 416898 589418 417134
rect 589502 416898 589738 417134
rect 589182 381218 589418 381454
rect 589502 381218 589738 381454
rect 589182 380898 589418 381134
rect 589502 380898 589738 381134
rect 589182 345218 589418 345454
rect 589502 345218 589738 345454
rect 589182 344898 589418 345134
rect 589502 344898 589738 345134
rect 589182 309218 589418 309454
rect 589502 309218 589738 309454
rect 589182 308898 589418 309134
rect 589502 308898 589738 309134
rect 589182 273218 589418 273454
rect 589502 273218 589738 273454
rect 589182 272898 589418 273134
rect 589502 272898 589738 273134
rect 589182 237218 589418 237454
rect 589502 237218 589738 237454
rect 589182 236898 589418 237134
rect 589502 236898 589738 237134
rect 589182 201218 589418 201454
rect 589502 201218 589738 201454
rect 589182 200898 589418 201134
rect 589502 200898 589738 201134
rect 589182 165218 589418 165454
rect 589502 165218 589738 165454
rect 589182 164898 589418 165134
rect 589502 164898 589738 165134
rect 589182 129218 589418 129454
rect 589502 129218 589738 129454
rect 589182 128898 589418 129134
rect 589502 128898 589738 129134
rect 589182 93218 589418 93454
rect 589502 93218 589738 93454
rect 589182 92898 589418 93134
rect 589502 92898 589738 93134
rect 589182 57218 589418 57454
rect 589502 57218 589738 57454
rect 589182 56898 589418 57134
rect 589502 56898 589738 57134
rect 589182 21218 589418 21454
rect 589502 21218 589738 21454
rect 589182 20898 589418 21134
rect 589502 20898 589738 21134
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 673718 590378 673954
rect 590462 673718 590698 673954
rect 590142 673398 590378 673634
rect 590462 673398 590698 673634
rect 590142 637718 590378 637954
rect 590462 637718 590698 637954
rect 590142 637398 590378 637634
rect 590462 637398 590698 637634
rect 590142 601718 590378 601954
rect 590462 601718 590698 601954
rect 590142 601398 590378 601634
rect 590462 601398 590698 601634
rect 590142 565718 590378 565954
rect 590462 565718 590698 565954
rect 590142 565398 590378 565634
rect 590462 565398 590698 565634
rect 590142 529718 590378 529954
rect 590462 529718 590698 529954
rect 590142 529398 590378 529634
rect 590462 529398 590698 529634
rect 590142 493718 590378 493954
rect 590462 493718 590698 493954
rect 590142 493398 590378 493634
rect 590462 493398 590698 493634
rect 590142 457718 590378 457954
rect 590462 457718 590698 457954
rect 590142 457398 590378 457634
rect 590462 457398 590698 457634
rect 590142 421718 590378 421954
rect 590462 421718 590698 421954
rect 590142 421398 590378 421634
rect 590462 421398 590698 421634
rect 590142 385718 590378 385954
rect 590462 385718 590698 385954
rect 590142 385398 590378 385634
rect 590462 385398 590698 385634
rect 590142 349718 590378 349954
rect 590462 349718 590698 349954
rect 590142 349398 590378 349634
rect 590462 349398 590698 349634
rect 590142 313718 590378 313954
rect 590462 313718 590698 313954
rect 590142 313398 590378 313634
rect 590462 313398 590698 313634
rect 590142 277718 590378 277954
rect 590462 277718 590698 277954
rect 590142 277398 590378 277634
rect 590462 277398 590698 277634
rect 590142 241718 590378 241954
rect 590462 241718 590698 241954
rect 590142 241398 590378 241634
rect 590462 241398 590698 241634
rect 590142 205718 590378 205954
rect 590462 205718 590698 205954
rect 590142 205398 590378 205634
rect 590462 205398 590698 205634
rect 590142 169718 590378 169954
rect 590462 169718 590698 169954
rect 590142 169398 590378 169634
rect 590462 169398 590698 169634
rect 590142 133718 590378 133954
rect 590462 133718 590698 133954
rect 590142 133398 590378 133634
rect 590462 133398 590698 133634
rect 590142 97718 590378 97954
rect 590462 97718 590698 97954
rect 590142 97398 590378 97634
rect 590462 97398 590698 97634
rect 590142 61718 590378 61954
rect 590462 61718 590698 61954
rect 590142 61398 590378 61634
rect 590462 61398 590698 61634
rect 590142 25718 590378 25954
rect 590462 25718 590698 25954
rect 590142 25398 590378 25634
rect 590462 25398 590698 25634
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 678218 591338 678454
rect 591422 678218 591658 678454
rect 591102 677898 591338 678134
rect 591422 677898 591658 678134
rect 591102 642218 591338 642454
rect 591422 642218 591658 642454
rect 591102 641898 591338 642134
rect 591422 641898 591658 642134
rect 591102 606218 591338 606454
rect 591422 606218 591658 606454
rect 591102 605898 591338 606134
rect 591422 605898 591658 606134
rect 591102 570218 591338 570454
rect 591422 570218 591658 570454
rect 591102 569898 591338 570134
rect 591422 569898 591658 570134
rect 591102 534218 591338 534454
rect 591422 534218 591658 534454
rect 591102 533898 591338 534134
rect 591422 533898 591658 534134
rect 591102 498218 591338 498454
rect 591422 498218 591658 498454
rect 591102 497898 591338 498134
rect 591422 497898 591658 498134
rect 591102 462218 591338 462454
rect 591422 462218 591658 462454
rect 591102 461898 591338 462134
rect 591422 461898 591658 462134
rect 591102 426218 591338 426454
rect 591422 426218 591658 426454
rect 591102 425898 591338 426134
rect 591422 425898 591658 426134
rect 591102 390218 591338 390454
rect 591422 390218 591658 390454
rect 591102 389898 591338 390134
rect 591422 389898 591658 390134
rect 591102 354218 591338 354454
rect 591422 354218 591658 354454
rect 591102 353898 591338 354134
rect 591422 353898 591658 354134
rect 591102 318218 591338 318454
rect 591422 318218 591658 318454
rect 591102 317898 591338 318134
rect 591422 317898 591658 318134
rect 591102 282218 591338 282454
rect 591422 282218 591658 282454
rect 591102 281898 591338 282134
rect 591422 281898 591658 282134
rect 591102 246218 591338 246454
rect 591422 246218 591658 246454
rect 591102 245898 591338 246134
rect 591422 245898 591658 246134
rect 591102 210218 591338 210454
rect 591422 210218 591658 210454
rect 591102 209898 591338 210134
rect 591422 209898 591658 210134
rect 591102 174218 591338 174454
rect 591422 174218 591658 174454
rect 591102 173898 591338 174134
rect 591422 173898 591658 174134
rect 591102 138218 591338 138454
rect 591422 138218 591658 138454
rect 591102 137898 591338 138134
rect 591422 137898 591658 138134
rect 591102 102218 591338 102454
rect 591422 102218 591658 102454
rect 591102 101898 591338 102134
rect 591422 101898 591658 102134
rect 591102 66218 591338 66454
rect 591422 66218 591658 66454
rect 591102 65898 591338 66134
rect 591422 65898 591658 66134
rect 591102 30218 591338 30454
rect 591422 30218 591658 30454
rect 591102 29898 591338 30134
rect 591422 29898 591658 30134
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 682718 592298 682954
rect 592382 682718 592618 682954
rect 592062 682398 592298 682634
rect 592382 682398 592618 682634
rect 592062 646718 592298 646954
rect 592382 646718 592618 646954
rect 592062 646398 592298 646634
rect 592382 646398 592618 646634
rect 592062 610718 592298 610954
rect 592382 610718 592618 610954
rect 592062 610398 592298 610634
rect 592382 610398 592618 610634
rect 592062 574718 592298 574954
rect 592382 574718 592618 574954
rect 592062 574398 592298 574634
rect 592382 574398 592618 574634
rect 592062 538718 592298 538954
rect 592382 538718 592618 538954
rect 592062 538398 592298 538634
rect 592382 538398 592618 538634
rect 592062 502718 592298 502954
rect 592382 502718 592618 502954
rect 592062 502398 592298 502634
rect 592382 502398 592618 502634
rect 592062 466718 592298 466954
rect 592382 466718 592618 466954
rect 592062 466398 592298 466634
rect 592382 466398 592618 466634
rect 592062 430718 592298 430954
rect 592382 430718 592618 430954
rect 592062 430398 592298 430634
rect 592382 430398 592618 430634
rect 592062 394718 592298 394954
rect 592382 394718 592618 394954
rect 592062 394398 592298 394634
rect 592382 394398 592618 394634
rect 592062 358718 592298 358954
rect 592382 358718 592618 358954
rect 592062 358398 592298 358634
rect 592382 358398 592618 358634
rect 592062 322718 592298 322954
rect 592382 322718 592618 322954
rect 592062 322398 592298 322634
rect 592382 322398 592618 322634
rect 592062 286718 592298 286954
rect 592382 286718 592618 286954
rect 592062 286398 592298 286634
rect 592382 286398 592618 286634
rect 592062 250718 592298 250954
rect 592382 250718 592618 250954
rect 592062 250398 592298 250634
rect 592382 250398 592618 250634
rect 592062 214718 592298 214954
rect 592382 214718 592618 214954
rect 592062 214398 592298 214634
rect 592382 214398 592618 214634
rect 592062 178718 592298 178954
rect 592382 178718 592618 178954
rect 592062 178398 592298 178634
rect 592382 178398 592618 178634
rect 592062 142718 592298 142954
rect 592382 142718 592618 142954
rect 592062 142398 592298 142634
rect 592382 142398 592618 142634
rect 592062 106718 592298 106954
rect 592382 106718 592618 106954
rect 592062 106398 592298 106634
rect 592382 106398 592618 106634
rect 592062 70718 592298 70954
rect 592382 70718 592618 70954
rect 592062 70398 592298 70634
rect 592382 70398 592618 70634
rect 592062 34718 592298 34954
rect 592382 34718 592618 34954
rect 592062 34398 592298 34634
rect 592382 34398 592618 34634
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 33326 711558
rect 33562 711322 33646 711558
rect 33882 711322 69326 711558
rect 69562 711322 69646 711558
rect 69882 711322 105326 711558
rect 105562 711322 105646 711558
rect 105882 711322 141326 711558
rect 141562 711322 141646 711558
rect 141882 711322 177326 711558
rect 177562 711322 177646 711558
rect 177882 711322 213326 711558
rect 213562 711322 213646 711558
rect 213882 711322 249326 711558
rect 249562 711322 249646 711558
rect 249882 711322 285326 711558
rect 285562 711322 285646 711558
rect 285882 711322 321326 711558
rect 321562 711322 321646 711558
rect 321882 711322 357326 711558
rect 357562 711322 357646 711558
rect 357882 711322 393326 711558
rect 393562 711322 393646 711558
rect 393882 711322 429326 711558
rect 429562 711322 429646 711558
rect 429882 711322 465326 711558
rect 465562 711322 465646 711558
rect 465882 711322 501326 711558
rect 501562 711322 501646 711558
rect 501882 711322 537326 711558
rect 537562 711322 537646 711558
rect 537882 711322 573326 711558
rect 573562 711322 573646 711558
rect 573882 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 33326 711238
rect 33562 711002 33646 711238
rect 33882 711002 69326 711238
rect 69562 711002 69646 711238
rect 69882 711002 105326 711238
rect 105562 711002 105646 711238
rect 105882 711002 141326 711238
rect 141562 711002 141646 711238
rect 141882 711002 177326 711238
rect 177562 711002 177646 711238
rect 177882 711002 213326 711238
rect 213562 711002 213646 711238
rect 213882 711002 249326 711238
rect 249562 711002 249646 711238
rect 249882 711002 285326 711238
rect 285562 711002 285646 711238
rect 285882 711002 321326 711238
rect 321562 711002 321646 711238
rect 321882 711002 357326 711238
rect 357562 711002 357646 711238
rect 357882 711002 393326 711238
rect 393562 711002 393646 711238
rect 393882 711002 429326 711238
rect 429562 711002 429646 711238
rect 429882 711002 465326 711238
rect 465562 711002 465646 711238
rect 465882 711002 501326 711238
rect 501562 711002 501646 711238
rect 501882 711002 537326 711238
rect 537562 711002 537646 711238
rect 537882 711002 573326 711238
rect 573562 711002 573646 711238
rect 573882 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 28826 710598
rect 29062 710362 29146 710598
rect 29382 710362 64826 710598
rect 65062 710362 65146 710598
rect 65382 710362 100826 710598
rect 101062 710362 101146 710598
rect 101382 710362 136826 710598
rect 137062 710362 137146 710598
rect 137382 710362 172826 710598
rect 173062 710362 173146 710598
rect 173382 710362 208826 710598
rect 209062 710362 209146 710598
rect 209382 710362 244826 710598
rect 245062 710362 245146 710598
rect 245382 710362 280826 710598
rect 281062 710362 281146 710598
rect 281382 710362 316826 710598
rect 317062 710362 317146 710598
rect 317382 710362 352826 710598
rect 353062 710362 353146 710598
rect 353382 710362 388826 710598
rect 389062 710362 389146 710598
rect 389382 710362 424826 710598
rect 425062 710362 425146 710598
rect 425382 710362 460826 710598
rect 461062 710362 461146 710598
rect 461382 710362 496826 710598
rect 497062 710362 497146 710598
rect 497382 710362 532826 710598
rect 533062 710362 533146 710598
rect 533382 710362 568826 710598
rect 569062 710362 569146 710598
rect 569382 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 28826 710278
rect 29062 710042 29146 710278
rect 29382 710042 64826 710278
rect 65062 710042 65146 710278
rect 65382 710042 100826 710278
rect 101062 710042 101146 710278
rect 101382 710042 136826 710278
rect 137062 710042 137146 710278
rect 137382 710042 172826 710278
rect 173062 710042 173146 710278
rect 173382 710042 208826 710278
rect 209062 710042 209146 710278
rect 209382 710042 244826 710278
rect 245062 710042 245146 710278
rect 245382 710042 280826 710278
rect 281062 710042 281146 710278
rect 281382 710042 316826 710278
rect 317062 710042 317146 710278
rect 317382 710042 352826 710278
rect 353062 710042 353146 710278
rect 353382 710042 388826 710278
rect 389062 710042 389146 710278
rect 389382 710042 424826 710278
rect 425062 710042 425146 710278
rect 425382 710042 460826 710278
rect 461062 710042 461146 710278
rect 461382 710042 496826 710278
rect 497062 710042 497146 710278
rect 497382 710042 532826 710278
rect 533062 710042 533146 710278
rect 533382 710042 568826 710278
rect 569062 710042 569146 710278
rect 569382 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 24326 709638
rect 24562 709402 24646 709638
rect 24882 709402 60326 709638
rect 60562 709402 60646 709638
rect 60882 709402 96326 709638
rect 96562 709402 96646 709638
rect 96882 709402 132326 709638
rect 132562 709402 132646 709638
rect 132882 709402 168326 709638
rect 168562 709402 168646 709638
rect 168882 709402 204326 709638
rect 204562 709402 204646 709638
rect 204882 709402 240326 709638
rect 240562 709402 240646 709638
rect 240882 709402 276326 709638
rect 276562 709402 276646 709638
rect 276882 709402 312326 709638
rect 312562 709402 312646 709638
rect 312882 709402 348326 709638
rect 348562 709402 348646 709638
rect 348882 709402 384326 709638
rect 384562 709402 384646 709638
rect 384882 709402 420326 709638
rect 420562 709402 420646 709638
rect 420882 709402 456326 709638
rect 456562 709402 456646 709638
rect 456882 709402 492326 709638
rect 492562 709402 492646 709638
rect 492882 709402 528326 709638
rect 528562 709402 528646 709638
rect 528882 709402 564326 709638
rect 564562 709402 564646 709638
rect 564882 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 24326 709318
rect 24562 709082 24646 709318
rect 24882 709082 60326 709318
rect 60562 709082 60646 709318
rect 60882 709082 96326 709318
rect 96562 709082 96646 709318
rect 96882 709082 132326 709318
rect 132562 709082 132646 709318
rect 132882 709082 168326 709318
rect 168562 709082 168646 709318
rect 168882 709082 204326 709318
rect 204562 709082 204646 709318
rect 204882 709082 240326 709318
rect 240562 709082 240646 709318
rect 240882 709082 276326 709318
rect 276562 709082 276646 709318
rect 276882 709082 312326 709318
rect 312562 709082 312646 709318
rect 312882 709082 348326 709318
rect 348562 709082 348646 709318
rect 348882 709082 384326 709318
rect 384562 709082 384646 709318
rect 384882 709082 420326 709318
rect 420562 709082 420646 709318
rect 420882 709082 456326 709318
rect 456562 709082 456646 709318
rect 456882 709082 492326 709318
rect 492562 709082 492646 709318
rect 492882 709082 528326 709318
rect 528562 709082 528646 709318
rect 528882 709082 564326 709318
rect 564562 709082 564646 709318
rect 564882 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 19826 708678
rect 20062 708442 20146 708678
rect 20382 708442 55826 708678
rect 56062 708442 56146 708678
rect 56382 708442 91826 708678
rect 92062 708442 92146 708678
rect 92382 708442 127826 708678
rect 128062 708442 128146 708678
rect 128382 708442 163826 708678
rect 164062 708442 164146 708678
rect 164382 708442 199826 708678
rect 200062 708442 200146 708678
rect 200382 708442 235826 708678
rect 236062 708442 236146 708678
rect 236382 708442 271826 708678
rect 272062 708442 272146 708678
rect 272382 708442 307826 708678
rect 308062 708442 308146 708678
rect 308382 708442 343826 708678
rect 344062 708442 344146 708678
rect 344382 708442 379826 708678
rect 380062 708442 380146 708678
rect 380382 708442 415826 708678
rect 416062 708442 416146 708678
rect 416382 708442 451826 708678
rect 452062 708442 452146 708678
rect 452382 708442 487826 708678
rect 488062 708442 488146 708678
rect 488382 708442 523826 708678
rect 524062 708442 524146 708678
rect 524382 708442 559826 708678
rect 560062 708442 560146 708678
rect 560382 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 19826 708358
rect 20062 708122 20146 708358
rect 20382 708122 55826 708358
rect 56062 708122 56146 708358
rect 56382 708122 91826 708358
rect 92062 708122 92146 708358
rect 92382 708122 127826 708358
rect 128062 708122 128146 708358
rect 128382 708122 163826 708358
rect 164062 708122 164146 708358
rect 164382 708122 199826 708358
rect 200062 708122 200146 708358
rect 200382 708122 235826 708358
rect 236062 708122 236146 708358
rect 236382 708122 271826 708358
rect 272062 708122 272146 708358
rect 272382 708122 307826 708358
rect 308062 708122 308146 708358
rect 308382 708122 343826 708358
rect 344062 708122 344146 708358
rect 344382 708122 379826 708358
rect 380062 708122 380146 708358
rect 380382 708122 415826 708358
rect 416062 708122 416146 708358
rect 416382 708122 451826 708358
rect 452062 708122 452146 708358
rect 452382 708122 487826 708358
rect 488062 708122 488146 708358
rect 488382 708122 523826 708358
rect 524062 708122 524146 708358
rect 524382 708122 559826 708358
rect 560062 708122 560146 708358
rect 560382 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 15326 707718
rect 15562 707482 15646 707718
rect 15882 707482 51326 707718
rect 51562 707482 51646 707718
rect 51882 707482 87326 707718
rect 87562 707482 87646 707718
rect 87882 707482 123326 707718
rect 123562 707482 123646 707718
rect 123882 707482 159326 707718
rect 159562 707482 159646 707718
rect 159882 707482 195326 707718
rect 195562 707482 195646 707718
rect 195882 707482 231326 707718
rect 231562 707482 231646 707718
rect 231882 707482 267326 707718
rect 267562 707482 267646 707718
rect 267882 707482 303326 707718
rect 303562 707482 303646 707718
rect 303882 707482 339326 707718
rect 339562 707482 339646 707718
rect 339882 707482 375326 707718
rect 375562 707482 375646 707718
rect 375882 707482 411326 707718
rect 411562 707482 411646 707718
rect 411882 707482 447326 707718
rect 447562 707482 447646 707718
rect 447882 707482 483326 707718
rect 483562 707482 483646 707718
rect 483882 707482 519326 707718
rect 519562 707482 519646 707718
rect 519882 707482 555326 707718
rect 555562 707482 555646 707718
rect 555882 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 15326 707398
rect 15562 707162 15646 707398
rect 15882 707162 51326 707398
rect 51562 707162 51646 707398
rect 51882 707162 87326 707398
rect 87562 707162 87646 707398
rect 87882 707162 123326 707398
rect 123562 707162 123646 707398
rect 123882 707162 159326 707398
rect 159562 707162 159646 707398
rect 159882 707162 195326 707398
rect 195562 707162 195646 707398
rect 195882 707162 231326 707398
rect 231562 707162 231646 707398
rect 231882 707162 267326 707398
rect 267562 707162 267646 707398
rect 267882 707162 303326 707398
rect 303562 707162 303646 707398
rect 303882 707162 339326 707398
rect 339562 707162 339646 707398
rect 339882 707162 375326 707398
rect 375562 707162 375646 707398
rect 375882 707162 411326 707398
rect 411562 707162 411646 707398
rect 411882 707162 447326 707398
rect 447562 707162 447646 707398
rect 447882 707162 483326 707398
rect 483562 707162 483646 707398
rect 483882 707162 519326 707398
rect 519562 707162 519646 707398
rect 519882 707162 555326 707398
rect 555562 707162 555646 707398
rect 555882 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 10826 706758
rect 11062 706522 11146 706758
rect 11382 706522 46826 706758
rect 47062 706522 47146 706758
rect 47382 706522 82826 706758
rect 83062 706522 83146 706758
rect 83382 706522 118826 706758
rect 119062 706522 119146 706758
rect 119382 706522 154826 706758
rect 155062 706522 155146 706758
rect 155382 706522 190826 706758
rect 191062 706522 191146 706758
rect 191382 706522 226826 706758
rect 227062 706522 227146 706758
rect 227382 706522 262826 706758
rect 263062 706522 263146 706758
rect 263382 706522 298826 706758
rect 299062 706522 299146 706758
rect 299382 706522 334826 706758
rect 335062 706522 335146 706758
rect 335382 706522 370826 706758
rect 371062 706522 371146 706758
rect 371382 706522 406826 706758
rect 407062 706522 407146 706758
rect 407382 706522 442826 706758
rect 443062 706522 443146 706758
rect 443382 706522 478826 706758
rect 479062 706522 479146 706758
rect 479382 706522 514826 706758
rect 515062 706522 515146 706758
rect 515382 706522 550826 706758
rect 551062 706522 551146 706758
rect 551382 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 10826 706438
rect 11062 706202 11146 706438
rect 11382 706202 46826 706438
rect 47062 706202 47146 706438
rect 47382 706202 82826 706438
rect 83062 706202 83146 706438
rect 83382 706202 118826 706438
rect 119062 706202 119146 706438
rect 119382 706202 154826 706438
rect 155062 706202 155146 706438
rect 155382 706202 190826 706438
rect 191062 706202 191146 706438
rect 191382 706202 226826 706438
rect 227062 706202 227146 706438
rect 227382 706202 262826 706438
rect 263062 706202 263146 706438
rect 263382 706202 298826 706438
rect 299062 706202 299146 706438
rect 299382 706202 334826 706438
rect 335062 706202 335146 706438
rect 335382 706202 370826 706438
rect 371062 706202 371146 706438
rect 371382 706202 406826 706438
rect 407062 706202 407146 706438
rect 407382 706202 442826 706438
rect 443062 706202 443146 706438
rect 443382 706202 478826 706438
rect 479062 706202 479146 706438
rect 479382 706202 514826 706438
rect 515062 706202 515146 706438
rect 515382 706202 550826 706438
rect 551062 706202 551146 706438
rect 551382 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 6326 705798
rect 6562 705562 6646 705798
rect 6882 705562 42326 705798
rect 42562 705562 42646 705798
rect 42882 705562 78326 705798
rect 78562 705562 78646 705798
rect 78882 705562 114326 705798
rect 114562 705562 114646 705798
rect 114882 705562 150326 705798
rect 150562 705562 150646 705798
rect 150882 705562 186326 705798
rect 186562 705562 186646 705798
rect 186882 705562 222326 705798
rect 222562 705562 222646 705798
rect 222882 705562 258326 705798
rect 258562 705562 258646 705798
rect 258882 705562 294326 705798
rect 294562 705562 294646 705798
rect 294882 705562 330326 705798
rect 330562 705562 330646 705798
rect 330882 705562 366326 705798
rect 366562 705562 366646 705798
rect 366882 705562 402326 705798
rect 402562 705562 402646 705798
rect 402882 705562 438326 705798
rect 438562 705562 438646 705798
rect 438882 705562 474326 705798
rect 474562 705562 474646 705798
rect 474882 705562 510326 705798
rect 510562 705562 510646 705798
rect 510882 705562 546326 705798
rect 546562 705562 546646 705798
rect 546882 705562 582326 705798
rect 582562 705562 582646 705798
rect 582882 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 6326 705478
rect 6562 705242 6646 705478
rect 6882 705242 42326 705478
rect 42562 705242 42646 705478
rect 42882 705242 78326 705478
rect 78562 705242 78646 705478
rect 78882 705242 114326 705478
rect 114562 705242 114646 705478
rect 114882 705242 150326 705478
rect 150562 705242 150646 705478
rect 150882 705242 186326 705478
rect 186562 705242 186646 705478
rect 186882 705242 222326 705478
rect 222562 705242 222646 705478
rect 222882 705242 258326 705478
rect 258562 705242 258646 705478
rect 258882 705242 294326 705478
rect 294562 705242 294646 705478
rect 294882 705242 330326 705478
rect 330562 705242 330646 705478
rect 330882 705242 366326 705478
rect 366562 705242 366646 705478
rect 366882 705242 402326 705478
rect 402562 705242 402646 705478
rect 402882 705242 438326 705478
rect 438562 705242 438646 705478
rect 438882 705242 474326 705478
rect 474562 705242 474646 705478
rect 474882 705242 510326 705478
rect 510562 705242 510646 705478
rect 510882 705242 546326 705478
rect 546562 705242 546646 705478
rect 546882 705242 582326 705478
rect 582562 705242 582646 705478
rect 582882 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 700954 592650 700986
rect -8726 700718 -4854 700954
rect -4618 700718 -4534 700954
rect -4298 700718 15326 700954
rect 15562 700718 15646 700954
rect 15882 700718 51326 700954
rect 51562 700718 51646 700954
rect 51882 700718 87326 700954
rect 87562 700718 87646 700954
rect 87882 700718 123326 700954
rect 123562 700718 123646 700954
rect 123882 700718 159326 700954
rect 159562 700718 159646 700954
rect 159882 700718 195326 700954
rect 195562 700718 195646 700954
rect 195882 700718 231326 700954
rect 231562 700718 231646 700954
rect 231882 700718 267326 700954
rect 267562 700718 267646 700954
rect 267882 700718 303326 700954
rect 303562 700718 303646 700954
rect 303882 700718 339326 700954
rect 339562 700718 339646 700954
rect 339882 700718 375326 700954
rect 375562 700718 375646 700954
rect 375882 700718 411326 700954
rect 411562 700718 411646 700954
rect 411882 700718 447326 700954
rect 447562 700718 447646 700954
rect 447882 700718 483326 700954
rect 483562 700718 483646 700954
rect 483882 700718 519326 700954
rect 519562 700718 519646 700954
rect 519882 700718 555326 700954
rect 555562 700718 555646 700954
rect 555882 700718 588222 700954
rect 588458 700718 588542 700954
rect 588778 700718 592650 700954
rect -8726 700634 592650 700718
rect -8726 700398 -4854 700634
rect -4618 700398 -4534 700634
rect -4298 700398 15326 700634
rect 15562 700398 15646 700634
rect 15882 700398 51326 700634
rect 51562 700398 51646 700634
rect 51882 700398 87326 700634
rect 87562 700398 87646 700634
rect 87882 700398 123326 700634
rect 123562 700398 123646 700634
rect 123882 700398 159326 700634
rect 159562 700398 159646 700634
rect 159882 700398 195326 700634
rect 195562 700398 195646 700634
rect 195882 700398 231326 700634
rect 231562 700398 231646 700634
rect 231882 700398 267326 700634
rect 267562 700398 267646 700634
rect 267882 700398 303326 700634
rect 303562 700398 303646 700634
rect 303882 700398 339326 700634
rect 339562 700398 339646 700634
rect 339882 700398 375326 700634
rect 375562 700398 375646 700634
rect 375882 700398 411326 700634
rect 411562 700398 411646 700634
rect 411882 700398 447326 700634
rect 447562 700398 447646 700634
rect 447882 700398 483326 700634
rect 483562 700398 483646 700634
rect 483882 700398 519326 700634
rect 519562 700398 519646 700634
rect 519882 700398 555326 700634
rect 555562 700398 555646 700634
rect 555882 700398 588222 700634
rect 588458 700398 588542 700634
rect 588778 700398 592650 700634
rect -8726 700366 592650 700398
rect -8726 696454 592650 696486
rect -8726 696218 -3894 696454
rect -3658 696218 -3574 696454
rect -3338 696218 10826 696454
rect 11062 696218 11146 696454
rect 11382 696218 46826 696454
rect 47062 696218 47146 696454
rect 47382 696218 82826 696454
rect 83062 696218 83146 696454
rect 83382 696218 118826 696454
rect 119062 696218 119146 696454
rect 119382 696218 154826 696454
rect 155062 696218 155146 696454
rect 155382 696218 190826 696454
rect 191062 696218 191146 696454
rect 191382 696218 226826 696454
rect 227062 696218 227146 696454
rect 227382 696218 262826 696454
rect 263062 696218 263146 696454
rect 263382 696218 298826 696454
rect 299062 696218 299146 696454
rect 299382 696218 334826 696454
rect 335062 696218 335146 696454
rect 335382 696218 370826 696454
rect 371062 696218 371146 696454
rect 371382 696218 406826 696454
rect 407062 696218 407146 696454
rect 407382 696218 442826 696454
rect 443062 696218 443146 696454
rect 443382 696218 478826 696454
rect 479062 696218 479146 696454
rect 479382 696218 514826 696454
rect 515062 696218 515146 696454
rect 515382 696218 550826 696454
rect 551062 696218 551146 696454
rect 551382 696218 587262 696454
rect 587498 696218 587582 696454
rect 587818 696218 592650 696454
rect -8726 696134 592650 696218
rect -8726 695898 -3894 696134
rect -3658 695898 -3574 696134
rect -3338 695898 10826 696134
rect 11062 695898 11146 696134
rect 11382 695898 46826 696134
rect 47062 695898 47146 696134
rect 47382 695898 82826 696134
rect 83062 695898 83146 696134
rect 83382 695898 118826 696134
rect 119062 695898 119146 696134
rect 119382 695898 154826 696134
rect 155062 695898 155146 696134
rect 155382 695898 190826 696134
rect 191062 695898 191146 696134
rect 191382 695898 226826 696134
rect 227062 695898 227146 696134
rect 227382 695898 262826 696134
rect 263062 695898 263146 696134
rect 263382 695898 298826 696134
rect 299062 695898 299146 696134
rect 299382 695898 334826 696134
rect 335062 695898 335146 696134
rect 335382 695898 370826 696134
rect 371062 695898 371146 696134
rect 371382 695898 406826 696134
rect 407062 695898 407146 696134
rect 407382 695898 442826 696134
rect 443062 695898 443146 696134
rect 443382 695898 478826 696134
rect 479062 695898 479146 696134
rect 479382 695898 514826 696134
rect 515062 695898 515146 696134
rect 515382 695898 550826 696134
rect 551062 695898 551146 696134
rect 551382 695898 587262 696134
rect 587498 695898 587582 696134
rect 587818 695898 592650 696134
rect -8726 695866 592650 695898
rect -8726 691954 592650 691986
rect -8726 691718 -2934 691954
rect -2698 691718 -2614 691954
rect -2378 691718 6326 691954
rect 6562 691718 6646 691954
rect 6882 691718 42326 691954
rect 42562 691718 42646 691954
rect 42882 691718 78326 691954
rect 78562 691718 78646 691954
rect 78882 691718 114326 691954
rect 114562 691718 114646 691954
rect 114882 691718 150326 691954
rect 150562 691718 150646 691954
rect 150882 691718 186326 691954
rect 186562 691718 186646 691954
rect 186882 691718 222326 691954
rect 222562 691718 222646 691954
rect 222882 691718 258326 691954
rect 258562 691718 258646 691954
rect 258882 691718 294326 691954
rect 294562 691718 294646 691954
rect 294882 691718 330326 691954
rect 330562 691718 330646 691954
rect 330882 691718 366326 691954
rect 366562 691718 366646 691954
rect 366882 691718 402326 691954
rect 402562 691718 402646 691954
rect 402882 691718 438326 691954
rect 438562 691718 438646 691954
rect 438882 691718 474326 691954
rect 474562 691718 474646 691954
rect 474882 691718 510326 691954
rect 510562 691718 510646 691954
rect 510882 691718 546326 691954
rect 546562 691718 546646 691954
rect 546882 691718 582326 691954
rect 582562 691718 582646 691954
rect 582882 691718 586302 691954
rect 586538 691718 586622 691954
rect 586858 691718 592650 691954
rect -8726 691634 592650 691718
rect -8726 691398 -2934 691634
rect -2698 691398 -2614 691634
rect -2378 691398 6326 691634
rect 6562 691398 6646 691634
rect 6882 691398 42326 691634
rect 42562 691398 42646 691634
rect 42882 691398 78326 691634
rect 78562 691398 78646 691634
rect 78882 691398 114326 691634
rect 114562 691398 114646 691634
rect 114882 691398 150326 691634
rect 150562 691398 150646 691634
rect 150882 691398 186326 691634
rect 186562 691398 186646 691634
rect 186882 691398 222326 691634
rect 222562 691398 222646 691634
rect 222882 691398 258326 691634
rect 258562 691398 258646 691634
rect 258882 691398 294326 691634
rect 294562 691398 294646 691634
rect 294882 691398 330326 691634
rect 330562 691398 330646 691634
rect 330882 691398 366326 691634
rect 366562 691398 366646 691634
rect 366882 691398 402326 691634
rect 402562 691398 402646 691634
rect 402882 691398 438326 691634
rect 438562 691398 438646 691634
rect 438882 691398 474326 691634
rect 474562 691398 474646 691634
rect 474882 691398 510326 691634
rect 510562 691398 510646 691634
rect 510882 691398 546326 691634
rect 546562 691398 546646 691634
rect 546882 691398 582326 691634
rect 582562 691398 582646 691634
rect 582882 691398 586302 691634
rect 586538 691398 586622 691634
rect 586858 691398 592650 691634
rect -8726 691366 592650 691398
rect -8726 687454 592650 687486
rect -8726 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 592650 687454
rect -8726 687134 592650 687218
rect -8726 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 592650 687134
rect -8726 686866 592650 686898
rect -8726 682954 592650 682986
rect -8726 682718 -8694 682954
rect -8458 682718 -8374 682954
rect -8138 682718 33326 682954
rect 33562 682718 33646 682954
rect 33882 682718 69326 682954
rect 69562 682718 69646 682954
rect 69882 682718 105326 682954
rect 105562 682718 105646 682954
rect 105882 682718 141326 682954
rect 141562 682718 141646 682954
rect 141882 682718 177326 682954
rect 177562 682718 177646 682954
rect 177882 682718 213326 682954
rect 213562 682718 213646 682954
rect 213882 682718 249326 682954
rect 249562 682718 249646 682954
rect 249882 682718 285326 682954
rect 285562 682718 285646 682954
rect 285882 682718 321326 682954
rect 321562 682718 321646 682954
rect 321882 682718 357326 682954
rect 357562 682718 357646 682954
rect 357882 682718 393326 682954
rect 393562 682718 393646 682954
rect 393882 682718 429326 682954
rect 429562 682718 429646 682954
rect 429882 682718 465326 682954
rect 465562 682718 465646 682954
rect 465882 682718 501326 682954
rect 501562 682718 501646 682954
rect 501882 682718 537326 682954
rect 537562 682718 537646 682954
rect 537882 682718 573326 682954
rect 573562 682718 573646 682954
rect 573882 682718 592062 682954
rect 592298 682718 592382 682954
rect 592618 682718 592650 682954
rect -8726 682634 592650 682718
rect -8726 682398 -8694 682634
rect -8458 682398 -8374 682634
rect -8138 682398 33326 682634
rect 33562 682398 33646 682634
rect 33882 682398 69326 682634
rect 69562 682398 69646 682634
rect 69882 682398 105326 682634
rect 105562 682398 105646 682634
rect 105882 682398 141326 682634
rect 141562 682398 141646 682634
rect 141882 682398 177326 682634
rect 177562 682398 177646 682634
rect 177882 682398 213326 682634
rect 213562 682398 213646 682634
rect 213882 682398 249326 682634
rect 249562 682398 249646 682634
rect 249882 682398 285326 682634
rect 285562 682398 285646 682634
rect 285882 682398 321326 682634
rect 321562 682398 321646 682634
rect 321882 682398 357326 682634
rect 357562 682398 357646 682634
rect 357882 682398 393326 682634
rect 393562 682398 393646 682634
rect 393882 682398 429326 682634
rect 429562 682398 429646 682634
rect 429882 682398 465326 682634
rect 465562 682398 465646 682634
rect 465882 682398 501326 682634
rect 501562 682398 501646 682634
rect 501882 682398 537326 682634
rect 537562 682398 537646 682634
rect 537882 682398 573326 682634
rect 573562 682398 573646 682634
rect 573882 682398 592062 682634
rect 592298 682398 592382 682634
rect 592618 682398 592650 682634
rect -8726 682366 592650 682398
rect -8726 678454 592650 678486
rect -8726 678218 -7734 678454
rect -7498 678218 -7414 678454
rect -7178 678218 28826 678454
rect 29062 678218 29146 678454
rect 29382 678218 64826 678454
rect 65062 678218 65146 678454
rect 65382 678218 100826 678454
rect 101062 678218 101146 678454
rect 101382 678218 136826 678454
rect 137062 678218 137146 678454
rect 137382 678218 172826 678454
rect 173062 678218 173146 678454
rect 173382 678218 208826 678454
rect 209062 678218 209146 678454
rect 209382 678218 244826 678454
rect 245062 678218 245146 678454
rect 245382 678218 280826 678454
rect 281062 678218 281146 678454
rect 281382 678218 316826 678454
rect 317062 678218 317146 678454
rect 317382 678218 352826 678454
rect 353062 678218 353146 678454
rect 353382 678218 388826 678454
rect 389062 678218 389146 678454
rect 389382 678218 424826 678454
rect 425062 678218 425146 678454
rect 425382 678218 460826 678454
rect 461062 678218 461146 678454
rect 461382 678218 496826 678454
rect 497062 678218 497146 678454
rect 497382 678218 532826 678454
rect 533062 678218 533146 678454
rect 533382 678218 568826 678454
rect 569062 678218 569146 678454
rect 569382 678218 591102 678454
rect 591338 678218 591422 678454
rect 591658 678218 592650 678454
rect -8726 678134 592650 678218
rect -8726 677898 -7734 678134
rect -7498 677898 -7414 678134
rect -7178 677898 28826 678134
rect 29062 677898 29146 678134
rect 29382 677898 64826 678134
rect 65062 677898 65146 678134
rect 65382 677898 100826 678134
rect 101062 677898 101146 678134
rect 101382 677898 136826 678134
rect 137062 677898 137146 678134
rect 137382 677898 172826 678134
rect 173062 677898 173146 678134
rect 173382 677898 208826 678134
rect 209062 677898 209146 678134
rect 209382 677898 244826 678134
rect 245062 677898 245146 678134
rect 245382 677898 280826 678134
rect 281062 677898 281146 678134
rect 281382 677898 316826 678134
rect 317062 677898 317146 678134
rect 317382 677898 352826 678134
rect 353062 677898 353146 678134
rect 353382 677898 388826 678134
rect 389062 677898 389146 678134
rect 389382 677898 424826 678134
rect 425062 677898 425146 678134
rect 425382 677898 460826 678134
rect 461062 677898 461146 678134
rect 461382 677898 496826 678134
rect 497062 677898 497146 678134
rect 497382 677898 532826 678134
rect 533062 677898 533146 678134
rect 533382 677898 568826 678134
rect 569062 677898 569146 678134
rect 569382 677898 591102 678134
rect 591338 677898 591422 678134
rect 591658 677898 592650 678134
rect -8726 677866 592650 677898
rect -8726 673954 592650 673986
rect -8726 673718 -6774 673954
rect -6538 673718 -6454 673954
rect -6218 673718 24326 673954
rect 24562 673718 24646 673954
rect 24882 673718 60326 673954
rect 60562 673718 60646 673954
rect 60882 673718 96326 673954
rect 96562 673718 96646 673954
rect 96882 673718 132326 673954
rect 132562 673718 132646 673954
rect 132882 673718 168326 673954
rect 168562 673718 168646 673954
rect 168882 673718 204326 673954
rect 204562 673718 204646 673954
rect 204882 673718 240326 673954
rect 240562 673718 240646 673954
rect 240882 673718 276326 673954
rect 276562 673718 276646 673954
rect 276882 673718 312326 673954
rect 312562 673718 312646 673954
rect 312882 673718 348326 673954
rect 348562 673718 348646 673954
rect 348882 673718 384326 673954
rect 384562 673718 384646 673954
rect 384882 673718 420326 673954
rect 420562 673718 420646 673954
rect 420882 673718 456326 673954
rect 456562 673718 456646 673954
rect 456882 673718 492326 673954
rect 492562 673718 492646 673954
rect 492882 673718 528326 673954
rect 528562 673718 528646 673954
rect 528882 673718 564326 673954
rect 564562 673718 564646 673954
rect 564882 673718 590142 673954
rect 590378 673718 590462 673954
rect 590698 673718 592650 673954
rect -8726 673634 592650 673718
rect -8726 673398 -6774 673634
rect -6538 673398 -6454 673634
rect -6218 673398 24326 673634
rect 24562 673398 24646 673634
rect 24882 673398 60326 673634
rect 60562 673398 60646 673634
rect 60882 673398 96326 673634
rect 96562 673398 96646 673634
rect 96882 673398 132326 673634
rect 132562 673398 132646 673634
rect 132882 673398 168326 673634
rect 168562 673398 168646 673634
rect 168882 673398 204326 673634
rect 204562 673398 204646 673634
rect 204882 673398 240326 673634
rect 240562 673398 240646 673634
rect 240882 673398 276326 673634
rect 276562 673398 276646 673634
rect 276882 673398 312326 673634
rect 312562 673398 312646 673634
rect 312882 673398 348326 673634
rect 348562 673398 348646 673634
rect 348882 673398 384326 673634
rect 384562 673398 384646 673634
rect 384882 673398 420326 673634
rect 420562 673398 420646 673634
rect 420882 673398 456326 673634
rect 456562 673398 456646 673634
rect 456882 673398 492326 673634
rect 492562 673398 492646 673634
rect 492882 673398 528326 673634
rect 528562 673398 528646 673634
rect 528882 673398 564326 673634
rect 564562 673398 564646 673634
rect 564882 673398 590142 673634
rect 590378 673398 590462 673634
rect 590698 673398 592650 673634
rect -8726 673366 592650 673398
rect -8726 669454 592650 669486
rect -8726 669218 -5814 669454
rect -5578 669218 -5494 669454
rect -5258 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 589182 669454
rect 589418 669218 589502 669454
rect 589738 669218 592650 669454
rect -8726 669134 592650 669218
rect -8726 668898 -5814 669134
rect -5578 668898 -5494 669134
rect -5258 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 589182 669134
rect 589418 668898 589502 669134
rect 589738 668898 592650 669134
rect -8726 668866 592650 668898
rect -8726 664954 592650 664986
rect -8726 664718 -4854 664954
rect -4618 664718 -4534 664954
rect -4298 664718 15326 664954
rect 15562 664718 15646 664954
rect 15882 664718 51326 664954
rect 51562 664718 51646 664954
rect 51882 664718 87326 664954
rect 87562 664718 87646 664954
rect 87882 664718 123326 664954
rect 123562 664718 123646 664954
rect 123882 664718 159326 664954
rect 159562 664718 159646 664954
rect 159882 664718 195326 664954
rect 195562 664718 195646 664954
rect 195882 664718 231326 664954
rect 231562 664718 231646 664954
rect 231882 664718 267326 664954
rect 267562 664718 267646 664954
rect 267882 664718 303326 664954
rect 303562 664718 303646 664954
rect 303882 664718 339326 664954
rect 339562 664718 339646 664954
rect 339882 664718 375326 664954
rect 375562 664718 375646 664954
rect 375882 664718 411326 664954
rect 411562 664718 411646 664954
rect 411882 664718 447326 664954
rect 447562 664718 447646 664954
rect 447882 664718 483326 664954
rect 483562 664718 483646 664954
rect 483882 664718 519326 664954
rect 519562 664718 519646 664954
rect 519882 664718 555326 664954
rect 555562 664718 555646 664954
rect 555882 664718 588222 664954
rect 588458 664718 588542 664954
rect 588778 664718 592650 664954
rect -8726 664634 592650 664718
rect -8726 664398 -4854 664634
rect -4618 664398 -4534 664634
rect -4298 664398 15326 664634
rect 15562 664398 15646 664634
rect 15882 664398 51326 664634
rect 51562 664398 51646 664634
rect 51882 664398 87326 664634
rect 87562 664398 87646 664634
rect 87882 664398 123326 664634
rect 123562 664398 123646 664634
rect 123882 664398 159326 664634
rect 159562 664398 159646 664634
rect 159882 664398 195326 664634
rect 195562 664398 195646 664634
rect 195882 664398 231326 664634
rect 231562 664398 231646 664634
rect 231882 664398 267326 664634
rect 267562 664398 267646 664634
rect 267882 664398 303326 664634
rect 303562 664398 303646 664634
rect 303882 664398 339326 664634
rect 339562 664398 339646 664634
rect 339882 664398 375326 664634
rect 375562 664398 375646 664634
rect 375882 664398 411326 664634
rect 411562 664398 411646 664634
rect 411882 664398 447326 664634
rect 447562 664398 447646 664634
rect 447882 664398 483326 664634
rect 483562 664398 483646 664634
rect 483882 664398 519326 664634
rect 519562 664398 519646 664634
rect 519882 664398 555326 664634
rect 555562 664398 555646 664634
rect 555882 664398 588222 664634
rect 588458 664398 588542 664634
rect 588778 664398 592650 664634
rect -8726 664366 592650 664398
rect -8726 660454 592650 660486
rect -8726 660218 -3894 660454
rect -3658 660218 -3574 660454
rect -3338 660218 10826 660454
rect 11062 660218 11146 660454
rect 11382 660218 46826 660454
rect 47062 660218 47146 660454
rect 47382 660218 82826 660454
rect 83062 660218 83146 660454
rect 83382 660218 118826 660454
rect 119062 660218 119146 660454
rect 119382 660218 154826 660454
rect 155062 660218 155146 660454
rect 155382 660218 190826 660454
rect 191062 660218 191146 660454
rect 191382 660218 226826 660454
rect 227062 660218 227146 660454
rect 227382 660218 262826 660454
rect 263062 660218 263146 660454
rect 263382 660218 298826 660454
rect 299062 660218 299146 660454
rect 299382 660218 334826 660454
rect 335062 660218 335146 660454
rect 335382 660218 370826 660454
rect 371062 660218 371146 660454
rect 371382 660218 406826 660454
rect 407062 660218 407146 660454
rect 407382 660218 442826 660454
rect 443062 660218 443146 660454
rect 443382 660218 478826 660454
rect 479062 660218 479146 660454
rect 479382 660218 514826 660454
rect 515062 660218 515146 660454
rect 515382 660218 550826 660454
rect 551062 660218 551146 660454
rect 551382 660218 587262 660454
rect 587498 660218 587582 660454
rect 587818 660218 592650 660454
rect -8726 660134 592650 660218
rect -8726 659898 -3894 660134
rect -3658 659898 -3574 660134
rect -3338 659898 10826 660134
rect 11062 659898 11146 660134
rect 11382 659898 46826 660134
rect 47062 659898 47146 660134
rect 47382 659898 82826 660134
rect 83062 659898 83146 660134
rect 83382 659898 118826 660134
rect 119062 659898 119146 660134
rect 119382 659898 154826 660134
rect 155062 659898 155146 660134
rect 155382 659898 190826 660134
rect 191062 659898 191146 660134
rect 191382 659898 226826 660134
rect 227062 659898 227146 660134
rect 227382 659898 262826 660134
rect 263062 659898 263146 660134
rect 263382 659898 298826 660134
rect 299062 659898 299146 660134
rect 299382 659898 334826 660134
rect 335062 659898 335146 660134
rect 335382 659898 370826 660134
rect 371062 659898 371146 660134
rect 371382 659898 406826 660134
rect 407062 659898 407146 660134
rect 407382 659898 442826 660134
rect 443062 659898 443146 660134
rect 443382 659898 478826 660134
rect 479062 659898 479146 660134
rect 479382 659898 514826 660134
rect 515062 659898 515146 660134
rect 515382 659898 550826 660134
rect 551062 659898 551146 660134
rect 551382 659898 587262 660134
rect 587498 659898 587582 660134
rect 587818 659898 592650 660134
rect -8726 659866 592650 659898
rect -8726 655954 592650 655986
rect -8726 655718 -2934 655954
rect -2698 655718 -2614 655954
rect -2378 655718 6326 655954
rect 6562 655718 6646 655954
rect 6882 655718 42326 655954
rect 42562 655718 42646 655954
rect 42882 655718 78326 655954
rect 78562 655718 78646 655954
rect 78882 655718 114326 655954
rect 114562 655718 114646 655954
rect 114882 655718 150326 655954
rect 150562 655718 150646 655954
rect 150882 655718 186326 655954
rect 186562 655718 186646 655954
rect 186882 655718 222326 655954
rect 222562 655718 222646 655954
rect 222882 655718 258326 655954
rect 258562 655718 258646 655954
rect 258882 655718 294326 655954
rect 294562 655718 294646 655954
rect 294882 655718 330326 655954
rect 330562 655718 330646 655954
rect 330882 655718 366326 655954
rect 366562 655718 366646 655954
rect 366882 655718 402326 655954
rect 402562 655718 402646 655954
rect 402882 655718 438326 655954
rect 438562 655718 438646 655954
rect 438882 655718 474326 655954
rect 474562 655718 474646 655954
rect 474882 655718 510326 655954
rect 510562 655718 510646 655954
rect 510882 655718 546326 655954
rect 546562 655718 546646 655954
rect 546882 655718 582326 655954
rect 582562 655718 582646 655954
rect 582882 655718 586302 655954
rect 586538 655718 586622 655954
rect 586858 655718 592650 655954
rect -8726 655634 592650 655718
rect -8726 655398 -2934 655634
rect -2698 655398 -2614 655634
rect -2378 655398 6326 655634
rect 6562 655398 6646 655634
rect 6882 655398 42326 655634
rect 42562 655398 42646 655634
rect 42882 655398 78326 655634
rect 78562 655398 78646 655634
rect 78882 655398 114326 655634
rect 114562 655398 114646 655634
rect 114882 655398 150326 655634
rect 150562 655398 150646 655634
rect 150882 655398 186326 655634
rect 186562 655398 186646 655634
rect 186882 655398 222326 655634
rect 222562 655398 222646 655634
rect 222882 655398 258326 655634
rect 258562 655398 258646 655634
rect 258882 655398 294326 655634
rect 294562 655398 294646 655634
rect 294882 655398 330326 655634
rect 330562 655398 330646 655634
rect 330882 655398 366326 655634
rect 366562 655398 366646 655634
rect 366882 655398 402326 655634
rect 402562 655398 402646 655634
rect 402882 655398 438326 655634
rect 438562 655398 438646 655634
rect 438882 655398 474326 655634
rect 474562 655398 474646 655634
rect 474882 655398 510326 655634
rect 510562 655398 510646 655634
rect 510882 655398 546326 655634
rect 546562 655398 546646 655634
rect 546882 655398 582326 655634
rect 582562 655398 582646 655634
rect 582882 655398 586302 655634
rect 586538 655398 586622 655634
rect 586858 655398 592650 655634
rect -8726 655366 592650 655398
rect -8726 651454 592650 651486
rect -8726 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 592650 651454
rect -8726 651134 592650 651218
rect -8726 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 592650 651134
rect -8726 650866 592650 650898
rect -8726 646954 592650 646986
rect -8726 646718 -8694 646954
rect -8458 646718 -8374 646954
rect -8138 646718 33326 646954
rect 33562 646718 33646 646954
rect 33882 646718 69326 646954
rect 69562 646718 69646 646954
rect 69882 646718 105326 646954
rect 105562 646718 105646 646954
rect 105882 646718 141326 646954
rect 141562 646718 141646 646954
rect 141882 646718 177326 646954
rect 177562 646718 177646 646954
rect 177882 646718 213326 646954
rect 213562 646718 213646 646954
rect 213882 646718 249326 646954
rect 249562 646718 249646 646954
rect 249882 646718 285326 646954
rect 285562 646718 285646 646954
rect 285882 646718 321326 646954
rect 321562 646718 321646 646954
rect 321882 646718 357326 646954
rect 357562 646718 357646 646954
rect 357882 646718 393326 646954
rect 393562 646718 393646 646954
rect 393882 646718 429326 646954
rect 429562 646718 429646 646954
rect 429882 646718 465326 646954
rect 465562 646718 465646 646954
rect 465882 646718 501326 646954
rect 501562 646718 501646 646954
rect 501882 646718 537326 646954
rect 537562 646718 537646 646954
rect 537882 646718 573326 646954
rect 573562 646718 573646 646954
rect 573882 646718 592062 646954
rect 592298 646718 592382 646954
rect 592618 646718 592650 646954
rect -8726 646634 592650 646718
rect -8726 646398 -8694 646634
rect -8458 646398 -8374 646634
rect -8138 646398 33326 646634
rect 33562 646398 33646 646634
rect 33882 646398 69326 646634
rect 69562 646398 69646 646634
rect 69882 646398 105326 646634
rect 105562 646398 105646 646634
rect 105882 646398 141326 646634
rect 141562 646398 141646 646634
rect 141882 646398 177326 646634
rect 177562 646398 177646 646634
rect 177882 646398 213326 646634
rect 213562 646398 213646 646634
rect 213882 646398 249326 646634
rect 249562 646398 249646 646634
rect 249882 646398 285326 646634
rect 285562 646398 285646 646634
rect 285882 646398 321326 646634
rect 321562 646398 321646 646634
rect 321882 646398 357326 646634
rect 357562 646398 357646 646634
rect 357882 646398 393326 646634
rect 393562 646398 393646 646634
rect 393882 646398 429326 646634
rect 429562 646398 429646 646634
rect 429882 646398 465326 646634
rect 465562 646398 465646 646634
rect 465882 646398 501326 646634
rect 501562 646398 501646 646634
rect 501882 646398 537326 646634
rect 537562 646398 537646 646634
rect 537882 646398 573326 646634
rect 573562 646398 573646 646634
rect 573882 646398 592062 646634
rect 592298 646398 592382 646634
rect 592618 646398 592650 646634
rect -8726 646366 592650 646398
rect -8726 642454 592650 642486
rect -8726 642218 -7734 642454
rect -7498 642218 -7414 642454
rect -7178 642218 28826 642454
rect 29062 642218 29146 642454
rect 29382 642218 64826 642454
rect 65062 642218 65146 642454
rect 65382 642218 100826 642454
rect 101062 642218 101146 642454
rect 101382 642218 136826 642454
rect 137062 642218 137146 642454
rect 137382 642218 172826 642454
rect 173062 642218 173146 642454
rect 173382 642218 208826 642454
rect 209062 642218 209146 642454
rect 209382 642218 244826 642454
rect 245062 642218 245146 642454
rect 245382 642218 280826 642454
rect 281062 642218 281146 642454
rect 281382 642218 316826 642454
rect 317062 642218 317146 642454
rect 317382 642218 352826 642454
rect 353062 642218 353146 642454
rect 353382 642218 388826 642454
rect 389062 642218 389146 642454
rect 389382 642218 424826 642454
rect 425062 642218 425146 642454
rect 425382 642218 460826 642454
rect 461062 642218 461146 642454
rect 461382 642218 496826 642454
rect 497062 642218 497146 642454
rect 497382 642218 532826 642454
rect 533062 642218 533146 642454
rect 533382 642218 568826 642454
rect 569062 642218 569146 642454
rect 569382 642218 591102 642454
rect 591338 642218 591422 642454
rect 591658 642218 592650 642454
rect -8726 642134 592650 642218
rect -8726 641898 -7734 642134
rect -7498 641898 -7414 642134
rect -7178 641898 28826 642134
rect 29062 641898 29146 642134
rect 29382 641898 64826 642134
rect 65062 641898 65146 642134
rect 65382 641898 100826 642134
rect 101062 641898 101146 642134
rect 101382 641898 136826 642134
rect 137062 641898 137146 642134
rect 137382 641898 172826 642134
rect 173062 641898 173146 642134
rect 173382 641898 208826 642134
rect 209062 641898 209146 642134
rect 209382 641898 244826 642134
rect 245062 641898 245146 642134
rect 245382 641898 280826 642134
rect 281062 641898 281146 642134
rect 281382 641898 316826 642134
rect 317062 641898 317146 642134
rect 317382 641898 352826 642134
rect 353062 641898 353146 642134
rect 353382 641898 388826 642134
rect 389062 641898 389146 642134
rect 389382 641898 424826 642134
rect 425062 641898 425146 642134
rect 425382 641898 460826 642134
rect 461062 641898 461146 642134
rect 461382 641898 496826 642134
rect 497062 641898 497146 642134
rect 497382 641898 532826 642134
rect 533062 641898 533146 642134
rect 533382 641898 568826 642134
rect 569062 641898 569146 642134
rect 569382 641898 591102 642134
rect 591338 641898 591422 642134
rect 591658 641898 592650 642134
rect -8726 641866 592650 641898
rect -8726 637954 592650 637986
rect -8726 637718 -6774 637954
rect -6538 637718 -6454 637954
rect -6218 637718 24326 637954
rect 24562 637718 24646 637954
rect 24882 637718 60326 637954
rect 60562 637718 60646 637954
rect 60882 637718 96326 637954
rect 96562 637718 96646 637954
rect 96882 637718 132326 637954
rect 132562 637718 132646 637954
rect 132882 637718 168326 637954
rect 168562 637718 168646 637954
rect 168882 637718 204326 637954
rect 204562 637718 204646 637954
rect 204882 637718 240326 637954
rect 240562 637718 240646 637954
rect 240882 637718 276326 637954
rect 276562 637718 276646 637954
rect 276882 637718 312326 637954
rect 312562 637718 312646 637954
rect 312882 637718 348326 637954
rect 348562 637718 348646 637954
rect 348882 637718 384326 637954
rect 384562 637718 384646 637954
rect 384882 637718 420326 637954
rect 420562 637718 420646 637954
rect 420882 637718 456326 637954
rect 456562 637718 456646 637954
rect 456882 637718 492326 637954
rect 492562 637718 492646 637954
rect 492882 637718 528326 637954
rect 528562 637718 528646 637954
rect 528882 637718 564326 637954
rect 564562 637718 564646 637954
rect 564882 637718 590142 637954
rect 590378 637718 590462 637954
rect 590698 637718 592650 637954
rect -8726 637634 592650 637718
rect -8726 637398 -6774 637634
rect -6538 637398 -6454 637634
rect -6218 637398 24326 637634
rect 24562 637398 24646 637634
rect 24882 637398 60326 637634
rect 60562 637398 60646 637634
rect 60882 637398 96326 637634
rect 96562 637398 96646 637634
rect 96882 637398 132326 637634
rect 132562 637398 132646 637634
rect 132882 637398 168326 637634
rect 168562 637398 168646 637634
rect 168882 637398 204326 637634
rect 204562 637398 204646 637634
rect 204882 637398 240326 637634
rect 240562 637398 240646 637634
rect 240882 637398 276326 637634
rect 276562 637398 276646 637634
rect 276882 637398 312326 637634
rect 312562 637398 312646 637634
rect 312882 637398 348326 637634
rect 348562 637398 348646 637634
rect 348882 637398 384326 637634
rect 384562 637398 384646 637634
rect 384882 637398 420326 637634
rect 420562 637398 420646 637634
rect 420882 637398 456326 637634
rect 456562 637398 456646 637634
rect 456882 637398 492326 637634
rect 492562 637398 492646 637634
rect 492882 637398 528326 637634
rect 528562 637398 528646 637634
rect 528882 637398 564326 637634
rect 564562 637398 564646 637634
rect 564882 637398 590142 637634
rect 590378 637398 590462 637634
rect 590698 637398 592650 637634
rect -8726 637366 592650 637398
rect -8726 633454 592650 633486
rect -8726 633218 -5814 633454
rect -5578 633218 -5494 633454
rect -5258 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 589182 633454
rect 589418 633218 589502 633454
rect 589738 633218 592650 633454
rect -8726 633134 592650 633218
rect -8726 632898 -5814 633134
rect -5578 632898 -5494 633134
rect -5258 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 589182 633134
rect 589418 632898 589502 633134
rect 589738 632898 592650 633134
rect -8726 632866 592650 632898
rect -8726 628954 592650 628986
rect -8726 628718 -4854 628954
rect -4618 628718 -4534 628954
rect -4298 628718 15326 628954
rect 15562 628718 15646 628954
rect 15882 628718 51326 628954
rect 51562 628718 51646 628954
rect 51882 628718 87326 628954
rect 87562 628718 87646 628954
rect 87882 628718 123326 628954
rect 123562 628718 123646 628954
rect 123882 628718 159326 628954
rect 159562 628718 159646 628954
rect 159882 628718 195326 628954
rect 195562 628718 195646 628954
rect 195882 628718 231326 628954
rect 231562 628718 231646 628954
rect 231882 628718 267326 628954
rect 267562 628718 267646 628954
rect 267882 628718 303326 628954
rect 303562 628718 303646 628954
rect 303882 628718 339326 628954
rect 339562 628718 339646 628954
rect 339882 628718 375326 628954
rect 375562 628718 375646 628954
rect 375882 628718 411326 628954
rect 411562 628718 411646 628954
rect 411882 628718 447326 628954
rect 447562 628718 447646 628954
rect 447882 628718 483326 628954
rect 483562 628718 483646 628954
rect 483882 628718 519326 628954
rect 519562 628718 519646 628954
rect 519882 628718 555326 628954
rect 555562 628718 555646 628954
rect 555882 628718 588222 628954
rect 588458 628718 588542 628954
rect 588778 628718 592650 628954
rect -8726 628634 592650 628718
rect -8726 628398 -4854 628634
rect -4618 628398 -4534 628634
rect -4298 628398 15326 628634
rect 15562 628398 15646 628634
rect 15882 628398 51326 628634
rect 51562 628398 51646 628634
rect 51882 628398 87326 628634
rect 87562 628398 87646 628634
rect 87882 628398 123326 628634
rect 123562 628398 123646 628634
rect 123882 628398 159326 628634
rect 159562 628398 159646 628634
rect 159882 628398 195326 628634
rect 195562 628398 195646 628634
rect 195882 628398 231326 628634
rect 231562 628398 231646 628634
rect 231882 628398 267326 628634
rect 267562 628398 267646 628634
rect 267882 628398 303326 628634
rect 303562 628398 303646 628634
rect 303882 628398 339326 628634
rect 339562 628398 339646 628634
rect 339882 628398 375326 628634
rect 375562 628398 375646 628634
rect 375882 628398 411326 628634
rect 411562 628398 411646 628634
rect 411882 628398 447326 628634
rect 447562 628398 447646 628634
rect 447882 628398 483326 628634
rect 483562 628398 483646 628634
rect 483882 628398 519326 628634
rect 519562 628398 519646 628634
rect 519882 628398 555326 628634
rect 555562 628398 555646 628634
rect 555882 628398 588222 628634
rect 588458 628398 588542 628634
rect 588778 628398 592650 628634
rect -8726 628366 592650 628398
rect -8726 624454 592650 624486
rect -8726 624218 -3894 624454
rect -3658 624218 -3574 624454
rect -3338 624218 10826 624454
rect 11062 624218 11146 624454
rect 11382 624218 46826 624454
rect 47062 624218 47146 624454
rect 47382 624218 82826 624454
rect 83062 624218 83146 624454
rect 83382 624218 118826 624454
rect 119062 624218 119146 624454
rect 119382 624218 154826 624454
rect 155062 624218 155146 624454
rect 155382 624218 190826 624454
rect 191062 624218 191146 624454
rect 191382 624218 226826 624454
rect 227062 624218 227146 624454
rect 227382 624218 262826 624454
rect 263062 624218 263146 624454
rect 263382 624218 298826 624454
rect 299062 624218 299146 624454
rect 299382 624218 334826 624454
rect 335062 624218 335146 624454
rect 335382 624218 370826 624454
rect 371062 624218 371146 624454
rect 371382 624218 406826 624454
rect 407062 624218 407146 624454
rect 407382 624218 442826 624454
rect 443062 624218 443146 624454
rect 443382 624218 478826 624454
rect 479062 624218 479146 624454
rect 479382 624218 514826 624454
rect 515062 624218 515146 624454
rect 515382 624218 550826 624454
rect 551062 624218 551146 624454
rect 551382 624218 587262 624454
rect 587498 624218 587582 624454
rect 587818 624218 592650 624454
rect -8726 624134 592650 624218
rect -8726 623898 -3894 624134
rect -3658 623898 -3574 624134
rect -3338 623898 10826 624134
rect 11062 623898 11146 624134
rect 11382 623898 46826 624134
rect 47062 623898 47146 624134
rect 47382 623898 82826 624134
rect 83062 623898 83146 624134
rect 83382 623898 118826 624134
rect 119062 623898 119146 624134
rect 119382 623898 154826 624134
rect 155062 623898 155146 624134
rect 155382 623898 190826 624134
rect 191062 623898 191146 624134
rect 191382 623898 226826 624134
rect 227062 623898 227146 624134
rect 227382 623898 262826 624134
rect 263062 623898 263146 624134
rect 263382 623898 298826 624134
rect 299062 623898 299146 624134
rect 299382 623898 334826 624134
rect 335062 623898 335146 624134
rect 335382 623898 370826 624134
rect 371062 623898 371146 624134
rect 371382 623898 406826 624134
rect 407062 623898 407146 624134
rect 407382 623898 442826 624134
rect 443062 623898 443146 624134
rect 443382 623898 478826 624134
rect 479062 623898 479146 624134
rect 479382 623898 514826 624134
rect 515062 623898 515146 624134
rect 515382 623898 550826 624134
rect 551062 623898 551146 624134
rect 551382 623898 587262 624134
rect 587498 623898 587582 624134
rect 587818 623898 592650 624134
rect -8726 623866 592650 623898
rect -8726 619954 592650 619986
rect -8726 619718 -2934 619954
rect -2698 619718 -2614 619954
rect -2378 619718 6326 619954
rect 6562 619718 6646 619954
rect 6882 619718 42326 619954
rect 42562 619718 42646 619954
rect 42882 619718 78326 619954
rect 78562 619718 78646 619954
rect 78882 619718 114326 619954
rect 114562 619718 114646 619954
rect 114882 619718 150326 619954
rect 150562 619718 150646 619954
rect 150882 619718 186326 619954
rect 186562 619718 186646 619954
rect 186882 619718 222326 619954
rect 222562 619718 222646 619954
rect 222882 619718 258326 619954
rect 258562 619718 258646 619954
rect 258882 619718 294326 619954
rect 294562 619718 294646 619954
rect 294882 619718 330326 619954
rect 330562 619718 330646 619954
rect 330882 619718 366326 619954
rect 366562 619718 366646 619954
rect 366882 619718 402326 619954
rect 402562 619718 402646 619954
rect 402882 619718 438326 619954
rect 438562 619718 438646 619954
rect 438882 619718 474326 619954
rect 474562 619718 474646 619954
rect 474882 619718 510326 619954
rect 510562 619718 510646 619954
rect 510882 619718 546326 619954
rect 546562 619718 546646 619954
rect 546882 619718 582326 619954
rect 582562 619718 582646 619954
rect 582882 619718 586302 619954
rect 586538 619718 586622 619954
rect 586858 619718 592650 619954
rect -8726 619634 592650 619718
rect -8726 619398 -2934 619634
rect -2698 619398 -2614 619634
rect -2378 619398 6326 619634
rect 6562 619398 6646 619634
rect 6882 619398 42326 619634
rect 42562 619398 42646 619634
rect 42882 619398 78326 619634
rect 78562 619398 78646 619634
rect 78882 619398 114326 619634
rect 114562 619398 114646 619634
rect 114882 619398 150326 619634
rect 150562 619398 150646 619634
rect 150882 619398 186326 619634
rect 186562 619398 186646 619634
rect 186882 619398 222326 619634
rect 222562 619398 222646 619634
rect 222882 619398 258326 619634
rect 258562 619398 258646 619634
rect 258882 619398 294326 619634
rect 294562 619398 294646 619634
rect 294882 619398 330326 619634
rect 330562 619398 330646 619634
rect 330882 619398 366326 619634
rect 366562 619398 366646 619634
rect 366882 619398 402326 619634
rect 402562 619398 402646 619634
rect 402882 619398 438326 619634
rect 438562 619398 438646 619634
rect 438882 619398 474326 619634
rect 474562 619398 474646 619634
rect 474882 619398 510326 619634
rect 510562 619398 510646 619634
rect 510882 619398 546326 619634
rect 546562 619398 546646 619634
rect 546882 619398 582326 619634
rect 582562 619398 582646 619634
rect 582882 619398 586302 619634
rect 586538 619398 586622 619634
rect 586858 619398 592650 619634
rect -8726 619366 592650 619398
rect -8726 615454 592650 615486
rect -8726 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 592650 615454
rect -8726 615134 592650 615218
rect -8726 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 592650 615134
rect -8726 614866 592650 614898
rect -8726 610954 592650 610986
rect -8726 610718 -8694 610954
rect -8458 610718 -8374 610954
rect -8138 610718 33326 610954
rect 33562 610718 33646 610954
rect 33882 610718 69326 610954
rect 69562 610718 69646 610954
rect 69882 610718 105326 610954
rect 105562 610718 105646 610954
rect 105882 610718 141326 610954
rect 141562 610718 141646 610954
rect 141882 610718 177326 610954
rect 177562 610718 177646 610954
rect 177882 610718 213326 610954
rect 213562 610718 213646 610954
rect 213882 610718 249326 610954
rect 249562 610718 249646 610954
rect 249882 610718 285326 610954
rect 285562 610718 285646 610954
rect 285882 610718 321326 610954
rect 321562 610718 321646 610954
rect 321882 610718 357326 610954
rect 357562 610718 357646 610954
rect 357882 610718 393326 610954
rect 393562 610718 393646 610954
rect 393882 610718 429326 610954
rect 429562 610718 429646 610954
rect 429882 610718 465326 610954
rect 465562 610718 465646 610954
rect 465882 610718 501326 610954
rect 501562 610718 501646 610954
rect 501882 610718 537326 610954
rect 537562 610718 537646 610954
rect 537882 610718 573326 610954
rect 573562 610718 573646 610954
rect 573882 610718 592062 610954
rect 592298 610718 592382 610954
rect 592618 610718 592650 610954
rect -8726 610634 592650 610718
rect -8726 610398 -8694 610634
rect -8458 610398 -8374 610634
rect -8138 610398 33326 610634
rect 33562 610398 33646 610634
rect 33882 610398 69326 610634
rect 69562 610398 69646 610634
rect 69882 610398 105326 610634
rect 105562 610398 105646 610634
rect 105882 610398 141326 610634
rect 141562 610398 141646 610634
rect 141882 610398 177326 610634
rect 177562 610398 177646 610634
rect 177882 610398 213326 610634
rect 213562 610398 213646 610634
rect 213882 610398 249326 610634
rect 249562 610398 249646 610634
rect 249882 610398 285326 610634
rect 285562 610398 285646 610634
rect 285882 610398 321326 610634
rect 321562 610398 321646 610634
rect 321882 610398 357326 610634
rect 357562 610398 357646 610634
rect 357882 610398 393326 610634
rect 393562 610398 393646 610634
rect 393882 610398 429326 610634
rect 429562 610398 429646 610634
rect 429882 610398 465326 610634
rect 465562 610398 465646 610634
rect 465882 610398 501326 610634
rect 501562 610398 501646 610634
rect 501882 610398 537326 610634
rect 537562 610398 537646 610634
rect 537882 610398 573326 610634
rect 573562 610398 573646 610634
rect 573882 610398 592062 610634
rect 592298 610398 592382 610634
rect 592618 610398 592650 610634
rect -8726 610366 592650 610398
rect -8726 606454 592650 606486
rect -8726 606218 -7734 606454
rect -7498 606218 -7414 606454
rect -7178 606218 28826 606454
rect 29062 606218 29146 606454
rect 29382 606218 64826 606454
rect 65062 606218 65146 606454
rect 65382 606218 100826 606454
rect 101062 606218 101146 606454
rect 101382 606218 136826 606454
rect 137062 606218 137146 606454
rect 137382 606218 172826 606454
rect 173062 606218 173146 606454
rect 173382 606218 208826 606454
rect 209062 606218 209146 606454
rect 209382 606218 244826 606454
rect 245062 606218 245146 606454
rect 245382 606218 280826 606454
rect 281062 606218 281146 606454
rect 281382 606218 316826 606454
rect 317062 606218 317146 606454
rect 317382 606218 352826 606454
rect 353062 606218 353146 606454
rect 353382 606218 388826 606454
rect 389062 606218 389146 606454
rect 389382 606218 424826 606454
rect 425062 606218 425146 606454
rect 425382 606218 460826 606454
rect 461062 606218 461146 606454
rect 461382 606218 496826 606454
rect 497062 606218 497146 606454
rect 497382 606218 532826 606454
rect 533062 606218 533146 606454
rect 533382 606218 568826 606454
rect 569062 606218 569146 606454
rect 569382 606218 591102 606454
rect 591338 606218 591422 606454
rect 591658 606218 592650 606454
rect -8726 606134 592650 606218
rect -8726 605898 -7734 606134
rect -7498 605898 -7414 606134
rect -7178 605898 28826 606134
rect 29062 605898 29146 606134
rect 29382 605898 64826 606134
rect 65062 605898 65146 606134
rect 65382 605898 100826 606134
rect 101062 605898 101146 606134
rect 101382 605898 136826 606134
rect 137062 605898 137146 606134
rect 137382 605898 172826 606134
rect 173062 605898 173146 606134
rect 173382 605898 208826 606134
rect 209062 605898 209146 606134
rect 209382 605898 244826 606134
rect 245062 605898 245146 606134
rect 245382 605898 280826 606134
rect 281062 605898 281146 606134
rect 281382 605898 316826 606134
rect 317062 605898 317146 606134
rect 317382 605898 352826 606134
rect 353062 605898 353146 606134
rect 353382 605898 388826 606134
rect 389062 605898 389146 606134
rect 389382 605898 424826 606134
rect 425062 605898 425146 606134
rect 425382 605898 460826 606134
rect 461062 605898 461146 606134
rect 461382 605898 496826 606134
rect 497062 605898 497146 606134
rect 497382 605898 532826 606134
rect 533062 605898 533146 606134
rect 533382 605898 568826 606134
rect 569062 605898 569146 606134
rect 569382 605898 591102 606134
rect 591338 605898 591422 606134
rect 591658 605898 592650 606134
rect -8726 605866 592650 605898
rect -8726 601954 592650 601986
rect -8726 601718 -6774 601954
rect -6538 601718 -6454 601954
rect -6218 601718 24326 601954
rect 24562 601718 24646 601954
rect 24882 601718 60326 601954
rect 60562 601718 60646 601954
rect 60882 601718 96326 601954
rect 96562 601718 96646 601954
rect 96882 601718 132326 601954
rect 132562 601718 132646 601954
rect 132882 601718 168326 601954
rect 168562 601718 168646 601954
rect 168882 601718 204326 601954
rect 204562 601718 204646 601954
rect 204882 601718 240326 601954
rect 240562 601718 240646 601954
rect 240882 601718 276326 601954
rect 276562 601718 276646 601954
rect 276882 601718 312326 601954
rect 312562 601718 312646 601954
rect 312882 601718 348326 601954
rect 348562 601718 348646 601954
rect 348882 601718 384326 601954
rect 384562 601718 384646 601954
rect 384882 601718 420326 601954
rect 420562 601718 420646 601954
rect 420882 601718 456326 601954
rect 456562 601718 456646 601954
rect 456882 601718 492326 601954
rect 492562 601718 492646 601954
rect 492882 601718 528326 601954
rect 528562 601718 528646 601954
rect 528882 601718 564326 601954
rect 564562 601718 564646 601954
rect 564882 601718 590142 601954
rect 590378 601718 590462 601954
rect 590698 601718 592650 601954
rect -8726 601634 592650 601718
rect -8726 601398 -6774 601634
rect -6538 601398 -6454 601634
rect -6218 601398 24326 601634
rect 24562 601398 24646 601634
rect 24882 601398 60326 601634
rect 60562 601398 60646 601634
rect 60882 601398 96326 601634
rect 96562 601398 96646 601634
rect 96882 601398 132326 601634
rect 132562 601398 132646 601634
rect 132882 601398 168326 601634
rect 168562 601398 168646 601634
rect 168882 601398 204326 601634
rect 204562 601398 204646 601634
rect 204882 601398 240326 601634
rect 240562 601398 240646 601634
rect 240882 601398 276326 601634
rect 276562 601398 276646 601634
rect 276882 601398 312326 601634
rect 312562 601398 312646 601634
rect 312882 601398 348326 601634
rect 348562 601398 348646 601634
rect 348882 601398 384326 601634
rect 384562 601398 384646 601634
rect 384882 601398 420326 601634
rect 420562 601398 420646 601634
rect 420882 601398 456326 601634
rect 456562 601398 456646 601634
rect 456882 601398 492326 601634
rect 492562 601398 492646 601634
rect 492882 601398 528326 601634
rect 528562 601398 528646 601634
rect 528882 601398 564326 601634
rect 564562 601398 564646 601634
rect 564882 601398 590142 601634
rect 590378 601398 590462 601634
rect 590698 601398 592650 601634
rect -8726 601366 592650 601398
rect -8726 597454 592650 597486
rect -8726 597218 -5814 597454
rect -5578 597218 -5494 597454
rect -5258 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 589182 597454
rect 589418 597218 589502 597454
rect 589738 597218 592650 597454
rect -8726 597134 592650 597218
rect -8726 596898 -5814 597134
rect -5578 596898 -5494 597134
rect -5258 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 589182 597134
rect 589418 596898 589502 597134
rect 589738 596898 592650 597134
rect -8726 596866 592650 596898
rect -8726 592954 592650 592986
rect -8726 592718 -4854 592954
rect -4618 592718 -4534 592954
rect -4298 592718 15326 592954
rect 15562 592718 15646 592954
rect 15882 592718 51326 592954
rect 51562 592718 51646 592954
rect 51882 592718 87326 592954
rect 87562 592718 87646 592954
rect 87882 592718 123326 592954
rect 123562 592718 123646 592954
rect 123882 592718 159326 592954
rect 159562 592718 159646 592954
rect 159882 592718 195326 592954
rect 195562 592718 195646 592954
rect 195882 592718 231326 592954
rect 231562 592718 231646 592954
rect 231882 592718 267326 592954
rect 267562 592718 267646 592954
rect 267882 592718 303326 592954
rect 303562 592718 303646 592954
rect 303882 592718 339326 592954
rect 339562 592718 339646 592954
rect 339882 592718 375326 592954
rect 375562 592718 375646 592954
rect 375882 592718 411326 592954
rect 411562 592718 411646 592954
rect 411882 592718 447326 592954
rect 447562 592718 447646 592954
rect 447882 592718 483326 592954
rect 483562 592718 483646 592954
rect 483882 592718 519326 592954
rect 519562 592718 519646 592954
rect 519882 592718 555326 592954
rect 555562 592718 555646 592954
rect 555882 592718 588222 592954
rect 588458 592718 588542 592954
rect 588778 592718 592650 592954
rect -8726 592634 592650 592718
rect -8726 592398 -4854 592634
rect -4618 592398 -4534 592634
rect -4298 592398 15326 592634
rect 15562 592398 15646 592634
rect 15882 592398 51326 592634
rect 51562 592398 51646 592634
rect 51882 592398 87326 592634
rect 87562 592398 87646 592634
rect 87882 592398 123326 592634
rect 123562 592398 123646 592634
rect 123882 592398 159326 592634
rect 159562 592398 159646 592634
rect 159882 592398 195326 592634
rect 195562 592398 195646 592634
rect 195882 592398 231326 592634
rect 231562 592398 231646 592634
rect 231882 592398 267326 592634
rect 267562 592398 267646 592634
rect 267882 592398 303326 592634
rect 303562 592398 303646 592634
rect 303882 592398 339326 592634
rect 339562 592398 339646 592634
rect 339882 592398 375326 592634
rect 375562 592398 375646 592634
rect 375882 592398 411326 592634
rect 411562 592398 411646 592634
rect 411882 592398 447326 592634
rect 447562 592398 447646 592634
rect 447882 592398 483326 592634
rect 483562 592398 483646 592634
rect 483882 592398 519326 592634
rect 519562 592398 519646 592634
rect 519882 592398 555326 592634
rect 555562 592398 555646 592634
rect 555882 592398 588222 592634
rect 588458 592398 588542 592634
rect 588778 592398 592650 592634
rect -8726 592366 592650 592398
rect -8726 588454 592650 588486
rect -8726 588218 -3894 588454
rect -3658 588218 -3574 588454
rect -3338 588218 10826 588454
rect 11062 588218 11146 588454
rect 11382 588218 46826 588454
rect 47062 588218 47146 588454
rect 47382 588218 82826 588454
rect 83062 588218 83146 588454
rect 83382 588218 226826 588454
rect 227062 588218 227146 588454
rect 227382 588218 262826 588454
rect 263062 588218 263146 588454
rect 263382 588218 298826 588454
rect 299062 588218 299146 588454
rect 299382 588218 334826 588454
rect 335062 588218 335146 588454
rect 335382 588218 370826 588454
rect 371062 588218 371146 588454
rect 371382 588218 478826 588454
rect 479062 588218 479146 588454
rect 479382 588218 514826 588454
rect 515062 588218 515146 588454
rect 515382 588218 550826 588454
rect 551062 588218 551146 588454
rect 551382 588218 587262 588454
rect 587498 588218 587582 588454
rect 587818 588218 592650 588454
rect -8726 588134 592650 588218
rect -8726 587898 -3894 588134
rect -3658 587898 -3574 588134
rect -3338 587898 10826 588134
rect 11062 587898 11146 588134
rect 11382 587898 46826 588134
rect 47062 587898 47146 588134
rect 47382 587898 82826 588134
rect 83062 587898 83146 588134
rect 83382 587898 226826 588134
rect 227062 587898 227146 588134
rect 227382 587898 262826 588134
rect 263062 587898 263146 588134
rect 263382 587898 298826 588134
rect 299062 587898 299146 588134
rect 299382 587898 334826 588134
rect 335062 587898 335146 588134
rect 335382 587898 370826 588134
rect 371062 587898 371146 588134
rect 371382 587898 478826 588134
rect 479062 587898 479146 588134
rect 479382 587898 514826 588134
rect 515062 587898 515146 588134
rect 515382 587898 550826 588134
rect 551062 587898 551146 588134
rect 551382 587898 587262 588134
rect 587498 587898 587582 588134
rect 587818 587898 592650 588134
rect -8726 587866 592650 587898
rect -8726 583954 592650 583986
rect -8726 583718 -2934 583954
rect -2698 583718 -2614 583954
rect -2378 583718 6326 583954
rect 6562 583718 6646 583954
rect 6882 583718 42326 583954
rect 42562 583718 42646 583954
rect 42882 583718 78326 583954
rect 78562 583718 78646 583954
rect 78882 583718 100328 583954
rect 100564 583718 190496 583954
rect 190732 583718 222326 583954
rect 222562 583718 222646 583954
rect 222882 583718 258326 583954
rect 258562 583718 258646 583954
rect 258882 583718 294326 583954
rect 294562 583718 294646 583954
rect 294882 583718 330326 583954
rect 330562 583718 330646 583954
rect 330882 583718 366326 583954
rect 366562 583718 366646 583954
rect 366882 583718 380328 583954
rect 380564 583718 470496 583954
rect 470732 583718 474326 583954
rect 474562 583718 474646 583954
rect 474882 583718 510326 583954
rect 510562 583718 510646 583954
rect 510882 583718 546326 583954
rect 546562 583718 546646 583954
rect 546882 583718 582326 583954
rect 582562 583718 582646 583954
rect 582882 583718 586302 583954
rect 586538 583718 586622 583954
rect 586858 583718 592650 583954
rect -8726 583634 592650 583718
rect -8726 583398 -2934 583634
rect -2698 583398 -2614 583634
rect -2378 583398 6326 583634
rect 6562 583398 6646 583634
rect 6882 583398 42326 583634
rect 42562 583398 42646 583634
rect 42882 583398 78326 583634
rect 78562 583398 78646 583634
rect 78882 583398 100328 583634
rect 100564 583398 190496 583634
rect 190732 583398 222326 583634
rect 222562 583398 222646 583634
rect 222882 583398 258326 583634
rect 258562 583398 258646 583634
rect 258882 583398 294326 583634
rect 294562 583398 294646 583634
rect 294882 583398 330326 583634
rect 330562 583398 330646 583634
rect 330882 583398 366326 583634
rect 366562 583398 366646 583634
rect 366882 583398 380328 583634
rect 380564 583398 470496 583634
rect 470732 583398 474326 583634
rect 474562 583398 474646 583634
rect 474882 583398 510326 583634
rect 510562 583398 510646 583634
rect 510882 583398 546326 583634
rect 546562 583398 546646 583634
rect 546882 583398 582326 583634
rect 582562 583398 582646 583634
rect 582882 583398 586302 583634
rect 586538 583398 586622 583634
rect 586858 583398 592650 583634
rect -8726 583366 592650 583398
rect -8726 579454 592650 579486
rect -8726 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 101008 579454
rect 101244 579218 189816 579454
rect 190052 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 381008 579454
rect 381244 579218 469816 579454
rect 470052 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 592650 579454
rect -8726 579134 592650 579218
rect -8726 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 101008 579134
rect 101244 578898 189816 579134
rect 190052 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 381008 579134
rect 381244 578898 469816 579134
rect 470052 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 592650 579134
rect -8726 578866 592650 578898
rect -8726 574954 592650 574986
rect -8726 574718 -8694 574954
rect -8458 574718 -8374 574954
rect -8138 574718 33326 574954
rect 33562 574718 33646 574954
rect 33882 574718 69326 574954
rect 69562 574718 69646 574954
rect 69882 574718 213326 574954
rect 213562 574718 213646 574954
rect 213882 574718 249326 574954
rect 249562 574718 249646 574954
rect 249882 574718 285326 574954
rect 285562 574718 285646 574954
rect 285882 574718 321326 574954
rect 321562 574718 321646 574954
rect 321882 574718 357326 574954
rect 357562 574718 357646 574954
rect 357882 574718 501326 574954
rect 501562 574718 501646 574954
rect 501882 574718 537326 574954
rect 537562 574718 537646 574954
rect 537882 574718 573326 574954
rect 573562 574718 573646 574954
rect 573882 574718 592062 574954
rect 592298 574718 592382 574954
rect 592618 574718 592650 574954
rect -8726 574634 592650 574718
rect -8726 574398 -8694 574634
rect -8458 574398 -8374 574634
rect -8138 574398 33326 574634
rect 33562 574398 33646 574634
rect 33882 574398 69326 574634
rect 69562 574398 69646 574634
rect 69882 574398 213326 574634
rect 213562 574398 213646 574634
rect 213882 574398 249326 574634
rect 249562 574398 249646 574634
rect 249882 574398 285326 574634
rect 285562 574398 285646 574634
rect 285882 574398 321326 574634
rect 321562 574398 321646 574634
rect 321882 574398 357326 574634
rect 357562 574398 357646 574634
rect 357882 574398 501326 574634
rect 501562 574398 501646 574634
rect 501882 574398 537326 574634
rect 537562 574398 537646 574634
rect 537882 574398 573326 574634
rect 573562 574398 573646 574634
rect 573882 574398 592062 574634
rect 592298 574398 592382 574634
rect 592618 574398 592650 574634
rect -8726 574366 592650 574398
rect -8726 570454 592650 570486
rect -8726 570218 -7734 570454
rect -7498 570218 -7414 570454
rect -7178 570218 28826 570454
rect 29062 570218 29146 570454
rect 29382 570218 64826 570454
rect 65062 570218 65146 570454
rect 65382 570218 208826 570454
rect 209062 570218 209146 570454
rect 209382 570218 244826 570454
rect 245062 570218 245146 570454
rect 245382 570218 280826 570454
rect 281062 570218 281146 570454
rect 281382 570218 316826 570454
rect 317062 570218 317146 570454
rect 317382 570218 352826 570454
rect 353062 570218 353146 570454
rect 353382 570218 496826 570454
rect 497062 570218 497146 570454
rect 497382 570218 532826 570454
rect 533062 570218 533146 570454
rect 533382 570218 568826 570454
rect 569062 570218 569146 570454
rect 569382 570218 591102 570454
rect 591338 570218 591422 570454
rect 591658 570218 592650 570454
rect -8726 570134 592650 570218
rect -8726 569898 -7734 570134
rect -7498 569898 -7414 570134
rect -7178 569898 28826 570134
rect 29062 569898 29146 570134
rect 29382 569898 64826 570134
rect 65062 569898 65146 570134
rect 65382 569898 208826 570134
rect 209062 569898 209146 570134
rect 209382 569898 244826 570134
rect 245062 569898 245146 570134
rect 245382 569898 280826 570134
rect 281062 569898 281146 570134
rect 281382 569898 316826 570134
rect 317062 569898 317146 570134
rect 317382 569898 352826 570134
rect 353062 569898 353146 570134
rect 353382 569898 496826 570134
rect 497062 569898 497146 570134
rect 497382 569898 532826 570134
rect 533062 569898 533146 570134
rect 533382 569898 568826 570134
rect 569062 569898 569146 570134
rect 569382 569898 591102 570134
rect 591338 569898 591422 570134
rect 591658 569898 592650 570134
rect -8726 569866 592650 569898
rect -8726 565954 592650 565986
rect -8726 565718 -6774 565954
rect -6538 565718 -6454 565954
rect -6218 565718 24326 565954
rect 24562 565718 24646 565954
rect 24882 565718 60326 565954
rect 60562 565718 60646 565954
rect 60882 565718 96326 565954
rect 96562 565718 96646 565954
rect 96882 565718 204326 565954
rect 204562 565718 204646 565954
rect 204882 565718 240326 565954
rect 240562 565718 240646 565954
rect 240882 565718 276326 565954
rect 276562 565718 276646 565954
rect 276882 565718 312326 565954
rect 312562 565718 312646 565954
rect 312882 565718 348326 565954
rect 348562 565718 348646 565954
rect 348882 565718 492326 565954
rect 492562 565718 492646 565954
rect 492882 565718 528326 565954
rect 528562 565718 528646 565954
rect 528882 565718 564326 565954
rect 564562 565718 564646 565954
rect 564882 565718 590142 565954
rect 590378 565718 590462 565954
rect 590698 565718 592650 565954
rect -8726 565634 592650 565718
rect -8726 565398 -6774 565634
rect -6538 565398 -6454 565634
rect -6218 565398 24326 565634
rect 24562 565398 24646 565634
rect 24882 565398 60326 565634
rect 60562 565398 60646 565634
rect 60882 565398 96326 565634
rect 96562 565398 96646 565634
rect 96882 565398 204326 565634
rect 204562 565398 204646 565634
rect 204882 565398 240326 565634
rect 240562 565398 240646 565634
rect 240882 565398 276326 565634
rect 276562 565398 276646 565634
rect 276882 565398 312326 565634
rect 312562 565398 312646 565634
rect 312882 565398 348326 565634
rect 348562 565398 348646 565634
rect 348882 565398 492326 565634
rect 492562 565398 492646 565634
rect 492882 565398 528326 565634
rect 528562 565398 528646 565634
rect 528882 565398 564326 565634
rect 564562 565398 564646 565634
rect 564882 565398 590142 565634
rect 590378 565398 590462 565634
rect 590698 565398 592650 565634
rect -8726 565366 592650 565398
rect -8726 561454 592650 561486
rect -8726 561218 -5814 561454
rect -5578 561218 -5494 561454
rect -5258 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 589182 561454
rect 589418 561218 589502 561454
rect 589738 561218 592650 561454
rect -8726 561134 592650 561218
rect -8726 560898 -5814 561134
rect -5578 560898 -5494 561134
rect -5258 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 589182 561134
rect 589418 560898 589502 561134
rect 589738 560898 592650 561134
rect -8726 560866 592650 560898
rect -8726 556954 592650 556986
rect -8726 556718 -4854 556954
rect -4618 556718 -4534 556954
rect -4298 556718 15326 556954
rect 15562 556718 15646 556954
rect 15882 556718 51326 556954
rect 51562 556718 51646 556954
rect 51882 556718 87326 556954
rect 87562 556718 87646 556954
rect 87882 556718 195326 556954
rect 195562 556718 195646 556954
rect 195882 556718 231326 556954
rect 231562 556718 231646 556954
rect 231882 556718 267326 556954
rect 267562 556718 267646 556954
rect 267882 556718 303326 556954
rect 303562 556718 303646 556954
rect 303882 556718 339326 556954
rect 339562 556718 339646 556954
rect 339882 556718 375326 556954
rect 375562 556718 375646 556954
rect 375882 556718 483326 556954
rect 483562 556718 483646 556954
rect 483882 556718 519326 556954
rect 519562 556718 519646 556954
rect 519882 556718 555326 556954
rect 555562 556718 555646 556954
rect 555882 556718 588222 556954
rect 588458 556718 588542 556954
rect 588778 556718 592650 556954
rect -8726 556634 592650 556718
rect -8726 556398 -4854 556634
rect -4618 556398 -4534 556634
rect -4298 556398 15326 556634
rect 15562 556398 15646 556634
rect 15882 556398 51326 556634
rect 51562 556398 51646 556634
rect 51882 556398 87326 556634
rect 87562 556398 87646 556634
rect 87882 556398 195326 556634
rect 195562 556398 195646 556634
rect 195882 556398 231326 556634
rect 231562 556398 231646 556634
rect 231882 556398 267326 556634
rect 267562 556398 267646 556634
rect 267882 556398 303326 556634
rect 303562 556398 303646 556634
rect 303882 556398 339326 556634
rect 339562 556398 339646 556634
rect 339882 556398 375326 556634
rect 375562 556398 375646 556634
rect 375882 556398 483326 556634
rect 483562 556398 483646 556634
rect 483882 556398 519326 556634
rect 519562 556398 519646 556634
rect 519882 556398 555326 556634
rect 555562 556398 555646 556634
rect 555882 556398 588222 556634
rect 588458 556398 588542 556634
rect 588778 556398 592650 556634
rect -8726 556366 592650 556398
rect -8726 552454 592650 552486
rect -8726 552218 -3894 552454
rect -3658 552218 -3574 552454
rect -3338 552218 10826 552454
rect 11062 552218 11146 552454
rect 11382 552218 46826 552454
rect 47062 552218 47146 552454
rect 47382 552218 82826 552454
rect 83062 552218 83146 552454
rect 83382 552218 226826 552454
rect 227062 552218 227146 552454
rect 227382 552218 262826 552454
rect 263062 552218 263146 552454
rect 263382 552218 298826 552454
rect 299062 552218 299146 552454
rect 299382 552218 334826 552454
rect 335062 552218 335146 552454
rect 335382 552218 370826 552454
rect 371062 552218 371146 552454
rect 371382 552218 478826 552454
rect 479062 552218 479146 552454
rect 479382 552218 514826 552454
rect 515062 552218 515146 552454
rect 515382 552218 550826 552454
rect 551062 552218 551146 552454
rect 551382 552218 587262 552454
rect 587498 552218 587582 552454
rect 587818 552218 592650 552454
rect -8726 552134 592650 552218
rect -8726 551898 -3894 552134
rect -3658 551898 -3574 552134
rect -3338 551898 10826 552134
rect 11062 551898 11146 552134
rect 11382 551898 46826 552134
rect 47062 551898 47146 552134
rect 47382 551898 82826 552134
rect 83062 551898 83146 552134
rect 83382 551898 226826 552134
rect 227062 551898 227146 552134
rect 227382 551898 262826 552134
rect 263062 551898 263146 552134
rect 263382 551898 298826 552134
rect 299062 551898 299146 552134
rect 299382 551898 334826 552134
rect 335062 551898 335146 552134
rect 335382 551898 370826 552134
rect 371062 551898 371146 552134
rect 371382 551898 478826 552134
rect 479062 551898 479146 552134
rect 479382 551898 514826 552134
rect 515062 551898 515146 552134
rect 515382 551898 550826 552134
rect 551062 551898 551146 552134
rect 551382 551898 587262 552134
rect 587498 551898 587582 552134
rect 587818 551898 592650 552134
rect -8726 551866 592650 551898
rect -8726 547954 592650 547986
rect -8726 547718 -2934 547954
rect -2698 547718 -2614 547954
rect -2378 547718 6326 547954
rect 6562 547718 6646 547954
rect 6882 547718 42326 547954
rect 42562 547718 42646 547954
rect 42882 547718 78326 547954
rect 78562 547718 78646 547954
rect 78882 547718 100328 547954
rect 100564 547718 190496 547954
rect 190732 547718 222326 547954
rect 222562 547718 222646 547954
rect 222882 547718 258326 547954
rect 258562 547718 258646 547954
rect 258882 547718 294326 547954
rect 294562 547718 294646 547954
rect 294882 547718 330326 547954
rect 330562 547718 330646 547954
rect 330882 547718 366326 547954
rect 366562 547718 366646 547954
rect 366882 547718 380328 547954
rect 380564 547718 470496 547954
rect 470732 547718 474326 547954
rect 474562 547718 474646 547954
rect 474882 547718 510326 547954
rect 510562 547718 510646 547954
rect 510882 547718 546326 547954
rect 546562 547718 546646 547954
rect 546882 547718 582326 547954
rect 582562 547718 582646 547954
rect 582882 547718 586302 547954
rect 586538 547718 586622 547954
rect 586858 547718 592650 547954
rect -8726 547634 592650 547718
rect -8726 547398 -2934 547634
rect -2698 547398 -2614 547634
rect -2378 547398 6326 547634
rect 6562 547398 6646 547634
rect 6882 547398 42326 547634
rect 42562 547398 42646 547634
rect 42882 547398 78326 547634
rect 78562 547398 78646 547634
rect 78882 547398 100328 547634
rect 100564 547398 190496 547634
rect 190732 547398 222326 547634
rect 222562 547398 222646 547634
rect 222882 547398 258326 547634
rect 258562 547398 258646 547634
rect 258882 547398 294326 547634
rect 294562 547398 294646 547634
rect 294882 547398 330326 547634
rect 330562 547398 330646 547634
rect 330882 547398 366326 547634
rect 366562 547398 366646 547634
rect 366882 547398 380328 547634
rect 380564 547398 470496 547634
rect 470732 547398 474326 547634
rect 474562 547398 474646 547634
rect 474882 547398 510326 547634
rect 510562 547398 510646 547634
rect 510882 547398 546326 547634
rect 546562 547398 546646 547634
rect 546882 547398 582326 547634
rect 582562 547398 582646 547634
rect 582882 547398 586302 547634
rect 586538 547398 586622 547634
rect 586858 547398 592650 547634
rect -8726 547366 592650 547398
rect -8726 543454 592650 543486
rect -8726 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 101008 543454
rect 101244 543218 189816 543454
rect 190052 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 381008 543454
rect 381244 543218 469816 543454
rect 470052 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 592650 543454
rect -8726 543134 592650 543218
rect -8726 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 101008 543134
rect 101244 542898 189816 543134
rect 190052 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 381008 543134
rect 381244 542898 469816 543134
rect 470052 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 592650 543134
rect -8726 542866 592650 542898
rect -8726 538954 592650 538986
rect -8726 538718 -8694 538954
rect -8458 538718 -8374 538954
rect -8138 538718 33326 538954
rect 33562 538718 33646 538954
rect 33882 538718 69326 538954
rect 69562 538718 69646 538954
rect 69882 538718 213326 538954
rect 213562 538718 213646 538954
rect 213882 538718 249326 538954
rect 249562 538718 249646 538954
rect 249882 538718 285326 538954
rect 285562 538718 285646 538954
rect 285882 538718 321326 538954
rect 321562 538718 321646 538954
rect 321882 538718 357326 538954
rect 357562 538718 357646 538954
rect 357882 538718 501326 538954
rect 501562 538718 501646 538954
rect 501882 538718 537326 538954
rect 537562 538718 537646 538954
rect 537882 538718 573326 538954
rect 573562 538718 573646 538954
rect 573882 538718 592062 538954
rect 592298 538718 592382 538954
rect 592618 538718 592650 538954
rect -8726 538634 592650 538718
rect -8726 538398 -8694 538634
rect -8458 538398 -8374 538634
rect -8138 538398 33326 538634
rect 33562 538398 33646 538634
rect 33882 538398 69326 538634
rect 69562 538398 69646 538634
rect 69882 538398 213326 538634
rect 213562 538398 213646 538634
rect 213882 538398 249326 538634
rect 249562 538398 249646 538634
rect 249882 538398 285326 538634
rect 285562 538398 285646 538634
rect 285882 538398 321326 538634
rect 321562 538398 321646 538634
rect 321882 538398 357326 538634
rect 357562 538398 357646 538634
rect 357882 538398 501326 538634
rect 501562 538398 501646 538634
rect 501882 538398 537326 538634
rect 537562 538398 537646 538634
rect 537882 538398 573326 538634
rect 573562 538398 573646 538634
rect 573882 538398 592062 538634
rect 592298 538398 592382 538634
rect 592618 538398 592650 538634
rect -8726 538366 592650 538398
rect -8726 534454 592650 534486
rect -8726 534218 -7734 534454
rect -7498 534218 -7414 534454
rect -7178 534218 28826 534454
rect 29062 534218 29146 534454
rect 29382 534218 64826 534454
rect 65062 534218 65146 534454
rect 65382 534218 208826 534454
rect 209062 534218 209146 534454
rect 209382 534218 244826 534454
rect 245062 534218 245146 534454
rect 245382 534218 280826 534454
rect 281062 534218 281146 534454
rect 281382 534218 316826 534454
rect 317062 534218 317146 534454
rect 317382 534218 352826 534454
rect 353062 534218 353146 534454
rect 353382 534218 496826 534454
rect 497062 534218 497146 534454
rect 497382 534218 532826 534454
rect 533062 534218 533146 534454
rect 533382 534218 568826 534454
rect 569062 534218 569146 534454
rect 569382 534218 591102 534454
rect 591338 534218 591422 534454
rect 591658 534218 592650 534454
rect -8726 534134 592650 534218
rect -8726 533898 -7734 534134
rect -7498 533898 -7414 534134
rect -7178 533898 28826 534134
rect 29062 533898 29146 534134
rect 29382 533898 64826 534134
rect 65062 533898 65146 534134
rect 65382 533898 208826 534134
rect 209062 533898 209146 534134
rect 209382 533898 244826 534134
rect 245062 533898 245146 534134
rect 245382 533898 280826 534134
rect 281062 533898 281146 534134
rect 281382 533898 316826 534134
rect 317062 533898 317146 534134
rect 317382 533898 352826 534134
rect 353062 533898 353146 534134
rect 353382 533898 496826 534134
rect 497062 533898 497146 534134
rect 497382 533898 532826 534134
rect 533062 533898 533146 534134
rect 533382 533898 568826 534134
rect 569062 533898 569146 534134
rect 569382 533898 591102 534134
rect 591338 533898 591422 534134
rect 591658 533898 592650 534134
rect -8726 533866 592650 533898
rect -8726 529954 592650 529986
rect -8726 529718 -6774 529954
rect -6538 529718 -6454 529954
rect -6218 529718 24326 529954
rect 24562 529718 24646 529954
rect 24882 529718 60326 529954
rect 60562 529718 60646 529954
rect 60882 529718 96326 529954
rect 96562 529718 96646 529954
rect 96882 529718 204326 529954
rect 204562 529718 204646 529954
rect 204882 529718 240326 529954
rect 240562 529718 240646 529954
rect 240882 529718 276326 529954
rect 276562 529718 276646 529954
rect 276882 529718 312326 529954
rect 312562 529718 312646 529954
rect 312882 529718 348326 529954
rect 348562 529718 348646 529954
rect 348882 529718 492326 529954
rect 492562 529718 492646 529954
rect 492882 529718 528326 529954
rect 528562 529718 528646 529954
rect 528882 529718 564326 529954
rect 564562 529718 564646 529954
rect 564882 529718 590142 529954
rect 590378 529718 590462 529954
rect 590698 529718 592650 529954
rect -8726 529634 592650 529718
rect -8726 529398 -6774 529634
rect -6538 529398 -6454 529634
rect -6218 529398 24326 529634
rect 24562 529398 24646 529634
rect 24882 529398 60326 529634
rect 60562 529398 60646 529634
rect 60882 529398 96326 529634
rect 96562 529398 96646 529634
rect 96882 529398 204326 529634
rect 204562 529398 204646 529634
rect 204882 529398 240326 529634
rect 240562 529398 240646 529634
rect 240882 529398 276326 529634
rect 276562 529398 276646 529634
rect 276882 529398 312326 529634
rect 312562 529398 312646 529634
rect 312882 529398 348326 529634
rect 348562 529398 348646 529634
rect 348882 529398 492326 529634
rect 492562 529398 492646 529634
rect 492882 529398 528326 529634
rect 528562 529398 528646 529634
rect 528882 529398 564326 529634
rect 564562 529398 564646 529634
rect 564882 529398 590142 529634
rect 590378 529398 590462 529634
rect 590698 529398 592650 529634
rect -8726 529366 592650 529398
rect -8726 525454 592650 525486
rect -8726 525218 -5814 525454
rect -5578 525218 -5494 525454
rect -5258 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 589182 525454
rect 589418 525218 589502 525454
rect 589738 525218 592650 525454
rect -8726 525134 592650 525218
rect -8726 524898 -5814 525134
rect -5578 524898 -5494 525134
rect -5258 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 589182 525134
rect 589418 524898 589502 525134
rect 589738 524898 592650 525134
rect -8726 524866 592650 524898
rect -8726 520954 592650 520986
rect -8726 520718 -4854 520954
rect -4618 520718 -4534 520954
rect -4298 520718 15326 520954
rect 15562 520718 15646 520954
rect 15882 520718 51326 520954
rect 51562 520718 51646 520954
rect 51882 520718 87326 520954
rect 87562 520718 87646 520954
rect 87882 520718 195326 520954
rect 195562 520718 195646 520954
rect 195882 520718 231326 520954
rect 231562 520718 231646 520954
rect 231882 520718 267326 520954
rect 267562 520718 267646 520954
rect 267882 520718 303326 520954
rect 303562 520718 303646 520954
rect 303882 520718 339326 520954
rect 339562 520718 339646 520954
rect 339882 520718 375326 520954
rect 375562 520718 375646 520954
rect 375882 520718 483326 520954
rect 483562 520718 483646 520954
rect 483882 520718 519326 520954
rect 519562 520718 519646 520954
rect 519882 520718 555326 520954
rect 555562 520718 555646 520954
rect 555882 520718 588222 520954
rect 588458 520718 588542 520954
rect 588778 520718 592650 520954
rect -8726 520634 592650 520718
rect -8726 520398 -4854 520634
rect -4618 520398 -4534 520634
rect -4298 520398 15326 520634
rect 15562 520398 15646 520634
rect 15882 520398 51326 520634
rect 51562 520398 51646 520634
rect 51882 520398 87326 520634
rect 87562 520398 87646 520634
rect 87882 520398 195326 520634
rect 195562 520398 195646 520634
rect 195882 520398 231326 520634
rect 231562 520398 231646 520634
rect 231882 520398 267326 520634
rect 267562 520398 267646 520634
rect 267882 520398 303326 520634
rect 303562 520398 303646 520634
rect 303882 520398 339326 520634
rect 339562 520398 339646 520634
rect 339882 520398 375326 520634
rect 375562 520398 375646 520634
rect 375882 520398 483326 520634
rect 483562 520398 483646 520634
rect 483882 520398 519326 520634
rect 519562 520398 519646 520634
rect 519882 520398 555326 520634
rect 555562 520398 555646 520634
rect 555882 520398 588222 520634
rect 588458 520398 588542 520634
rect 588778 520398 592650 520634
rect -8726 520366 592650 520398
rect -8726 516454 592650 516486
rect -8726 516218 -3894 516454
rect -3658 516218 -3574 516454
rect -3338 516218 10826 516454
rect 11062 516218 11146 516454
rect 11382 516218 46826 516454
rect 47062 516218 47146 516454
rect 47382 516218 82826 516454
rect 83062 516218 83146 516454
rect 83382 516218 226826 516454
rect 227062 516218 227146 516454
rect 227382 516218 262826 516454
rect 263062 516218 263146 516454
rect 263382 516218 298826 516454
rect 299062 516218 299146 516454
rect 299382 516218 334826 516454
rect 335062 516218 335146 516454
rect 335382 516218 370826 516454
rect 371062 516218 371146 516454
rect 371382 516218 478826 516454
rect 479062 516218 479146 516454
rect 479382 516218 514826 516454
rect 515062 516218 515146 516454
rect 515382 516218 550826 516454
rect 551062 516218 551146 516454
rect 551382 516218 587262 516454
rect 587498 516218 587582 516454
rect 587818 516218 592650 516454
rect -8726 516134 592650 516218
rect -8726 515898 -3894 516134
rect -3658 515898 -3574 516134
rect -3338 515898 10826 516134
rect 11062 515898 11146 516134
rect 11382 515898 46826 516134
rect 47062 515898 47146 516134
rect 47382 515898 82826 516134
rect 83062 515898 83146 516134
rect 83382 515898 226826 516134
rect 227062 515898 227146 516134
rect 227382 515898 262826 516134
rect 263062 515898 263146 516134
rect 263382 515898 298826 516134
rect 299062 515898 299146 516134
rect 299382 515898 334826 516134
rect 335062 515898 335146 516134
rect 335382 515898 370826 516134
rect 371062 515898 371146 516134
rect 371382 515898 478826 516134
rect 479062 515898 479146 516134
rect 479382 515898 514826 516134
rect 515062 515898 515146 516134
rect 515382 515898 550826 516134
rect 551062 515898 551146 516134
rect 551382 515898 587262 516134
rect 587498 515898 587582 516134
rect 587818 515898 592650 516134
rect -8726 515866 592650 515898
rect -8726 511954 592650 511986
rect -8726 511718 -2934 511954
rect -2698 511718 -2614 511954
rect -2378 511718 6326 511954
rect 6562 511718 6646 511954
rect 6882 511718 42326 511954
rect 42562 511718 42646 511954
rect 42882 511718 78326 511954
rect 78562 511718 78646 511954
rect 78882 511718 100328 511954
rect 100564 511718 190496 511954
rect 190732 511718 222326 511954
rect 222562 511718 222646 511954
rect 222882 511718 258326 511954
rect 258562 511718 258646 511954
rect 258882 511718 294326 511954
rect 294562 511718 294646 511954
rect 294882 511718 330326 511954
rect 330562 511718 330646 511954
rect 330882 511718 366326 511954
rect 366562 511718 366646 511954
rect 366882 511718 380328 511954
rect 380564 511718 470496 511954
rect 470732 511718 474326 511954
rect 474562 511718 474646 511954
rect 474882 511718 510326 511954
rect 510562 511718 510646 511954
rect 510882 511718 546326 511954
rect 546562 511718 546646 511954
rect 546882 511718 582326 511954
rect 582562 511718 582646 511954
rect 582882 511718 586302 511954
rect 586538 511718 586622 511954
rect 586858 511718 592650 511954
rect -8726 511634 592650 511718
rect -8726 511398 -2934 511634
rect -2698 511398 -2614 511634
rect -2378 511398 6326 511634
rect 6562 511398 6646 511634
rect 6882 511398 42326 511634
rect 42562 511398 42646 511634
rect 42882 511398 78326 511634
rect 78562 511398 78646 511634
rect 78882 511398 100328 511634
rect 100564 511398 190496 511634
rect 190732 511398 222326 511634
rect 222562 511398 222646 511634
rect 222882 511398 258326 511634
rect 258562 511398 258646 511634
rect 258882 511398 294326 511634
rect 294562 511398 294646 511634
rect 294882 511398 330326 511634
rect 330562 511398 330646 511634
rect 330882 511398 366326 511634
rect 366562 511398 366646 511634
rect 366882 511398 380328 511634
rect 380564 511398 470496 511634
rect 470732 511398 474326 511634
rect 474562 511398 474646 511634
rect 474882 511398 510326 511634
rect 510562 511398 510646 511634
rect 510882 511398 546326 511634
rect 546562 511398 546646 511634
rect 546882 511398 582326 511634
rect 582562 511398 582646 511634
rect 582882 511398 586302 511634
rect 586538 511398 586622 511634
rect 586858 511398 592650 511634
rect -8726 511366 592650 511398
rect -8726 507454 592650 507486
rect -8726 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 101008 507454
rect 101244 507218 189816 507454
rect 190052 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 381008 507454
rect 381244 507218 469816 507454
rect 470052 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 592650 507454
rect -8726 507134 592650 507218
rect -8726 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 101008 507134
rect 101244 506898 189816 507134
rect 190052 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 381008 507134
rect 381244 506898 469816 507134
rect 470052 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 592650 507134
rect -8726 506866 592650 506898
rect -8726 502954 592650 502986
rect -8726 502718 -8694 502954
rect -8458 502718 -8374 502954
rect -8138 502718 33326 502954
rect 33562 502718 33646 502954
rect 33882 502718 69326 502954
rect 69562 502718 69646 502954
rect 69882 502718 213326 502954
rect 213562 502718 213646 502954
rect 213882 502718 249326 502954
rect 249562 502718 249646 502954
rect 249882 502718 285326 502954
rect 285562 502718 285646 502954
rect 285882 502718 321326 502954
rect 321562 502718 321646 502954
rect 321882 502718 357326 502954
rect 357562 502718 357646 502954
rect 357882 502718 501326 502954
rect 501562 502718 501646 502954
rect 501882 502718 537326 502954
rect 537562 502718 537646 502954
rect 537882 502718 573326 502954
rect 573562 502718 573646 502954
rect 573882 502718 592062 502954
rect 592298 502718 592382 502954
rect 592618 502718 592650 502954
rect -8726 502634 592650 502718
rect -8726 502398 -8694 502634
rect -8458 502398 -8374 502634
rect -8138 502398 33326 502634
rect 33562 502398 33646 502634
rect 33882 502398 69326 502634
rect 69562 502398 69646 502634
rect 69882 502398 213326 502634
rect 213562 502398 213646 502634
rect 213882 502398 249326 502634
rect 249562 502398 249646 502634
rect 249882 502398 285326 502634
rect 285562 502398 285646 502634
rect 285882 502398 321326 502634
rect 321562 502398 321646 502634
rect 321882 502398 357326 502634
rect 357562 502398 357646 502634
rect 357882 502398 501326 502634
rect 501562 502398 501646 502634
rect 501882 502398 537326 502634
rect 537562 502398 537646 502634
rect 537882 502398 573326 502634
rect 573562 502398 573646 502634
rect 573882 502398 592062 502634
rect 592298 502398 592382 502634
rect 592618 502398 592650 502634
rect -8726 502366 592650 502398
rect -8726 498454 592650 498486
rect -8726 498218 -7734 498454
rect -7498 498218 -7414 498454
rect -7178 498218 28826 498454
rect 29062 498218 29146 498454
rect 29382 498218 64826 498454
rect 65062 498218 65146 498454
rect 65382 498218 208826 498454
rect 209062 498218 209146 498454
rect 209382 498218 244826 498454
rect 245062 498218 245146 498454
rect 245382 498218 280826 498454
rect 281062 498218 281146 498454
rect 281382 498218 316826 498454
rect 317062 498218 317146 498454
rect 317382 498218 352826 498454
rect 353062 498218 353146 498454
rect 353382 498218 496826 498454
rect 497062 498218 497146 498454
rect 497382 498218 532826 498454
rect 533062 498218 533146 498454
rect 533382 498218 568826 498454
rect 569062 498218 569146 498454
rect 569382 498218 591102 498454
rect 591338 498218 591422 498454
rect 591658 498218 592650 498454
rect -8726 498134 592650 498218
rect -8726 497898 -7734 498134
rect -7498 497898 -7414 498134
rect -7178 497898 28826 498134
rect 29062 497898 29146 498134
rect 29382 497898 64826 498134
rect 65062 497898 65146 498134
rect 65382 497898 208826 498134
rect 209062 497898 209146 498134
rect 209382 497898 244826 498134
rect 245062 497898 245146 498134
rect 245382 497898 280826 498134
rect 281062 497898 281146 498134
rect 281382 497898 316826 498134
rect 317062 497898 317146 498134
rect 317382 497898 352826 498134
rect 353062 497898 353146 498134
rect 353382 497898 496826 498134
rect 497062 497898 497146 498134
rect 497382 497898 532826 498134
rect 533062 497898 533146 498134
rect 533382 497898 568826 498134
rect 569062 497898 569146 498134
rect 569382 497898 591102 498134
rect 591338 497898 591422 498134
rect 591658 497898 592650 498134
rect -8726 497866 592650 497898
rect -8726 493954 592650 493986
rect -8726 493718 -6774 493954
rect -6538 493718 -6454 493954
rect -6218 493718 24326 493954
rect 24562 493718 24646 493954
rect 24882 493718 60326 493954
rect 60562 493718 60646 493954
rect 60882 493718 96326 493954
rect 96562 493718 96646 493954
rect 96882 493718 132326 493954
rect 132562 493718 132646 493954
rect 132882 493718 168326 493954
rect 168562 493718 168646 493954
rect 168882 493718 204326 493954
rect 204562 493718 204646 493954
rect 204882 493718 240326 493954
rect 240562 493718 240646 493954
rect 240882 493718 276326 493954
rect 276562 493718 276646 493954
rect 276882 493718 312326 493954
rect 312562 493718 312646 493954
rect 312882 493718 348326 493954
rect 348562 493718 348646 493954
rect 348882 493718 384326 493954
rect 384562 493718 384646 493954
rect 384882 493718 420326 493954
rect 420562 493718 420646 493954
rect 420882 493718 456326 493954
rect 456562 493718 456646 493954
rect 456882 493718 492326 493954
rect 492562 493718 492646 493954
rect 492882 493718 528326 493954
rect 528562 493718 528646 493954
rect 528882 493718 564326 493954
rect 564562 493718 564646 493954
rect 564882 493718 590142 493954
rect 590378 493718 590462 493954
rect 590698 493718 592650 493954
rect -8726 493634 592650 493718
rect -8726 493398 -6774 493634
rect -6538 493398 -6454 493634
rect -6218 493398 24326 493634
rect 24562 493398 24646 493634
rect 24882 493398 60326 493634
rect 60562 493398 60646 493634
rect 60882 493398 96326 493634
rect 96562 493398 96646 493634
rect 96882 493398 132326 493634
rect 132562 493398 132646 493634
rect 132882 493398 168326 493634
rect 168562 493398 168646 493634
rect 168882 493398 204326 493634
rect 204562 493398 204646 493634
rect 204882 493398 240326 493634
rect 240562 493398 240646 493634
rect 240882 493398 276326 493634
rect 276562 493398 276646 493634
rect 276882 493398 312326 493634
rect 312562 493398 312646 493634
rect 312882 493398 348326 493634
rect 348562 493398 348646 493634
rect 348882 493398 384326 493634
rect 384562 493398 384646 493634
rect 384882 493398 420326 493634
rect 420562 493398 420646 493634
rect 420882 493398 456326 493634
rect 456562 493398 456646 493634
rect 456882 493398 492326 493634
rect 492562 493398 492646 493634
rect 492882 493398 528326 493634
rect 528562 493398 528646 493634
rect 528882 493398 564326 493634
rect 564562 493398 564646 493634
rect 564882 493398 590142 493634
rect 590378 493398 590462 493634
rect 590698 493398 592650 493634
rect -8726 493366 592650 493398
rect -8726 489454 592650 489486
rect -8726 489218 -5814 489454
rect -5578 489218 -5494 489454
rect -5258 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 589182 489454
rect 589418 489218 589502 489454
rect 589738 489218 592650 489454
rect -8726 489134 592650 489218
rect -8726 488898 -5814 489134
rect -5578 488898 -5494 489134
rect -5258 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 589182 489134
rect 589418 488898 589502 489134
rect 589738 488898 592650 489134
rect -8726 488866 592650 488898
rect -8726 484954 592650 484986
rect -8726 484718 -4854 484954
rect -4618 484718 -4534 484954
rect -4298 484718 15326 484954
rect 15562 484718 15646 484954
rect 15882 484718 51326 484954
rect 51562 484718 51646 484954
rect 51882 484718 87326 484954
rect 87562 484718 87646 484954
rect 87882 484718 123326 484954
rect 123562 484718 123646 484954
rect 123882 484718 159326 484954
rect 159562 484718 159646 484954
rect 159882 484718 195326 484954
rect 195562 484718 195646 484954
rect 195882 484718 231326 484954
rect 231562 484718 231646 484954
rect 231882 484718 267326 484954
rect 267562 484718 267646 484954
rect 267882 484718 303326 484954
rect 303562 484718 303646 484954
rect 303882 484718 339326 484954
rect 339562 484718 339646 484954
rect 339882 484718 375326 484954
rect 375562 484718 375646 484954
rect 375882 484718 411326 484954
rect 411562 484718 411646 484954
rect 411882 484718 447326 484954
rect 447562 484718 447646 484954
rect 447882 484718 483326 484954
rect 483562 484718 483646 484954
rect 483882 484718 519326 484954
rect 519562 484718 519646 484954
rect 519882 484718 555326 484954
rect 555562 484718 555646 484954
rect 555882 484718 588222 484954
rect 588458 484718 588542 484954
rect 588778 484718 592650 484954
rect -8726 484634 592650 484718
rect -8726 484398 -4854 484634
rect -4618 484398 -4534 484634
rect -4298 484398 15326 484634
rect 15562 484398 15646 484634
rect 15882 484398 51326 484634
rect 51562 484398 51646 484634
rect 51882 484398 87326 484634
rect 87562 484398 87646 484634
rect 87882 484398 123326 484634
rect 123562 484398 123646 484634
rect 123882 484398 159326 484634
rect 159562 484398 159646 484634
rect 159882 484398 195326 484634
rect 195562 484398 195646 484634
rect 195882 484398 231326 484634
rect 231562 484398 231646 484634
rect 231882 484398 267326 484634
rect 267562 484398 267646 484634
rect 267882 484398 303326 484634
rect 303562 484398 303646 484634
rect 303882 484398 339326 484634
rect 339562 484398 339646 484634
rect 339882 484398 375326 484634
rect 375562 484398 375646 484634
rect 375882 484398 411326 484634
rect 411562 484398 411646 484634
rect 411882 484398 447326 484634
rect 447562 484398 447646 484634
rect 447882 484398 483326 484634
rect 483562 484398 483646 484634
rect 483882 484398 519326 484634
rect 519562 484398 519646 484634
rect 519882 484398 555326 484634
rect 555562 484398 555646 484634
rect 555882 484398 588222 484634
rect 588458 484398 588542 484634
rect 588778 484398 592650 484634
rect -8726 484366 592650 484398
rect -8726 480454 592650 480486
rect -8726 480218 -3894 480454
rect -3658 480218 -3574 480454
rect -3338 480218 10826 480454
rect 11062 480218 11146 480454
rect 11382 480218 46826 480454
rect 47062 480218 47146 480454
rect 47382 480218 82826 480454
rect 83062 480218 83146 480454
rect 83382 480218 118826 480454
rect 119062 480218 119146 480454
rect 119382 480218 154826 480454
rect 155062 480218 155146 480454
rect 155382 480218 190826 480454
rect 191062 480218 191146 480454
rect 191382 480218 226826 480454
rect 227062 480218 227146 480454
rect 227382 480218 262826 480454
rect 263062 480218 263146 480454
rect 263382 480218 298826 480454
rect 299062 480218 299146 480454
rect 299382 480218 334826 480454
rect 335062 480218 335146 480454
rect 335382 480218 370826 480454
rect 371062 480218 371146 480454
rect 371382 480218 406826 480454
rect 407062 480218 407146 480454
rect 407382 480218 442826 480454
rect 443062 480218 443146 480454
rect 443382 480218 478826 480454
rect 479062 480218 479146 480454
rect 479382 480218 514826 480454
rect 515062 480218 515146 480454
rect 515382 480218 550826 480454
rect 551062 480218 551146 480454
rect 551382 480218 587262 480454
rect 587498 480218 587582 480454
rect 587818 480218 592650 480454
rect -8726 480134 592650 480218
rect -8726 479898 -3894 480134
rect -3658 479898 -3574 480134
rect -3338 479898 10826 480134
rect 11062 479898 11146 480134
rect 11382 479898 46826 480134
rect 47062 479898 47146 480134
rect 47382 479898 82826 480134
rect 83062 479898 83146 480134
rect 83382 479898 118826 480134
rect 119062 479898 119146 480134
rect 119382 479898 154826 480134
rect 155062 479898 155146 480134
rect 155382 479898 190826 480134
rect 191062 479898 191146 480134
rect 191382 479898 226826 480134
rect 227062 479898 227146 480134
rect 227382 479898 262826 480134
rect 263062 479898 263146 480134
rect 263382 479898 298826 480134
rect 299062 479898 299146 480134
rect 299382 479898 334826 480134
rect 335062 479898 335146 480134
rect 335382 479898 370826 480134
rect 371062 479898 371146 480134
rect 371382 479898 406826 480134
rect 407062 479898 407146 480134
rect 407382 479898 442826 480134
rect 443062 479898 443146 480134
rect 443382 479898 478826 480134
rect 479062 479898 479146 480134
rect 479382 479898 514826 480134
rect 515062 479898 515146 480134
rect 515382 479898 550826 480134
rect 551062 479898 551146 480134
rect 551382 479898 587262 480134
rect 587498 479898 587582 480134
rect 587818 479898 592650 480134
rect -8726 479866 592650 479898
rect -8726 475954 592650 475986
rect -8726 475718 -2934 475954
rect -2698 475718 -2614 475954
rect -2378 475718 6326 475954
rect 6562 475718 6646 475954
rect 6882 475718 42326 475954
rect 42562 475718 42646 475954
rect 42882 475718 78326 475954
rect 78562 475718 78646 475954
rect 78882 475718 114326 475954
rect 114562 475718 114646 475954
rect 114882 475718 150326 475954
rect 150562 475718 150646 475954
rect 150882 475718 186326 475954
rect 186562 475718 186646 475954
rect 186882 475718 222326 475954
rect 222562 475718 222646 475954
rect 222882 475718 258326 475954
rect 258562 475718 258646 475954
rect 258882 475718 294326 475954
rect 294562 475718 294646 475954
rect 294882 475718 330326 475954
rect 330562 475718 330646 475954
rect 330882 475718 366326 475954
rect 366562 475718 366646 475954
rect 366882 475718 402326 475954
rect 402562 475718 402646 475954
rect 402882 475718 438326 475954
rect 438562 475718 438646 475954
rect 438882 475718 474326 475954
rect 474562 475718 474646 475954
rect 474882 475718 510326 475954
rect 510562 475718 510646 475954
rect 510882 475718 546326 475954
rect 546562 475718 546646 475954
rect 546882 475718 582326 475954
rect 582562 475718 582646 475954
rect 582882 475718 586302 475954
rect 586538 475718 586622 475954
rect 586858 475718 592650 475954
rect -8726 475634 592650 475718
rect -8726 475398 -2934 475634
rect -2698 475398 -2614 475634
rect -2378 475398 6326 475634
rect 6562 475398 6646 475634
rect 6882 475398 42326 475634
rect 42562 475398 42646 475634
rect 42882 475398 78326 475634
rect 78562 475398 78646 475634
rect 78882 475398 114326 475634
rect 114562 475398 114646 475634
rect 114882 475398 150326 475634
rect 150562 475398 150646 475634
rect 150882 475398 186326 475634
rect 186562 475398 186646 475634
rect 186882 475398 222326 475634
rect 222562 475398 222646 475634
rect 222882 475398 258326 475634
rect 258562 475398 258646 475634
rect 258882 475398 294326 475634
rect 294562 475398 294646 475634
rect 294882 475398 330326 475634
rect 330562 475398 330646 475634
rect 330882 475398 366326 475634
rect 366562 475398 366646 475634
rect 366882 475398 402326 475634
rect 402562 475398 402646 475634
rect 402882 475398 438326 475634
rect 438562 475398 438646 475634
rect 438882 475398 474326 475634
rect 474562 475398 474646 475634
rect 474882 475398 510326 475634
rect 510562 475398 510646 475634
rect 510882 475398 546326 475634
rect 546562 475398 546646 475634
rect 546882 475398 582326 475634
rect 582562 475398 582646 475634
rect 582882 475398 586302 475634
rect 586538 475398 586622 475634
rect 586858 475398 592650 475634
rect -8726 475366 592650 475398
rect -8726 471454 592650 471486
rect -8726 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 592650 471454
rect -8726 471134 592650 471218
rect -8726 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 592650 471134
rect -8726 470866 592650 470898
rect -8726 466954 592650 466986
rect -8726 466718 -8694 466954
rect -8458 466718 -8374 466954
rect -8138 466718 33326 466954
rect 33562 466718 33646 466954
rect 33882 466718 69326 466954
rect 69562 466718 69646 466954
rect 69882 466718 105326 466954
rect 105562 466718 105646 466954
rect 105882 466718 141326 466954
rect 141562 466718 141646 466954
rect 141882 466718 177326 466954
rect 177562 466718 177646 466954
rect 177882 466718 213326 466954
rect 213562 466718 213646 466954
rect 213882 466718 249326 466954
rect 249562 466718 249646 466954
rect 249882 466718 285326 466954
rect 285562 466718 285646 466954
rect 285882 466718 321326 466954
rect 321562 466718 321646 466954
rect 321882 466718 357326 466954
rect 357562 466718 357646 466954
rect 357882 466718 393326 466954
rect 393562 466718 393646 466954
rect 393882 466718 429326 466954
rect 429562 466718 429646 466954
rect 429882 466718 465326 466954
rect 465562 466718 465646 466954
rect 465882 466718 501326 466954
rect 501562 466718 501646 466954
rect 501882 466718 537326 466954
rect 537562 466718 537646 466954
rect 537882 466718 573326 466954
rect 573562 466718 573646 466954
rect 573882 466718 592062 466954
rect 592298 466718 592382 466954
rect 592618 466718 592650 466954
rect -8726 466634 592650 466718
rect -8726 466398 -8694 466634
rect -8458 466398 -8374 466634
rect -8138 466398 33326 466634
rect 33562 466398 33646 466634
rect 33882 466398 69326 466634
rect 69562 466398 69646 466634
rect 69882 466398 105326 466634
rect 105562 466398 105646 466634
rect 105882 466398 141326 466634
rect 141562 466398 141646 466634
rect 141882 466398 177326 466634
rect 177562 466398 177646 466634
rect 177882 466398 213326 466634
rect 213562 466398 213646 466634
rect 213882 466398 249326 466634
rect 249562 466398 249646 466634
rect 249882 466398 285326 466634
rect 285562 466398 285646 466634
rect 285882 466398 321326 466634
rect 321562 466398 321646 466634
rect 321882 466398 357326 466634
rect 357562 466398 357646 466634
rect 357882 466398 393326 466634
rect 393562 466398 393646 466634
rect 393882 466398 429326 466634
rect 429562 466398 429646 466634
rect 429882 466398 465326 466634
rect 465562 466398 465646 466634
rect 465882 466398 501326 466634
rect 501562 466398 501646 466634
rect 501882 466398 537326 466634
rect 537562 466398 537646 466634
rect 537882 466398 573326 466634
rect 573562 466398 573646 466634
rect 573882 466398 592062 466634
rect 592298 466398 592382 466634
rect 592618 466398 592650 466634
rect -8726 466366 592650 466398
rect -8726 462454 592650 462486
rect -8726 462218 -7734 462454
rect -7498 462218 -7414 462454
rect -7178 462218 28826 462454
rect 29062 462218 29146 462454
rect 29382 462218 64826 462454
rect 65062 462218 65146 462454
rect 65382 462218 100826 462454
rect 101062 462218 101146 462454
rect 101382 462218 136826 462454
rect 137062 462218 137146 462454
rect 137382 462218 172826 462454
rect 173062 462218 173146 462454
rect 173382 462218 208826 462454
rect 209062 462218 209146 462454
rect 209382 462218 244826 462454
rect 245062 462218 245146 462454
rect 245382 462218 280826 462454
rect 281062 462218 281146 462454
rect 281382 462218 316826 462454
rect 317062 462218 317146 462454
rect 317382 462218 352826 462454
rect 353062 462218 353146 462454
rect 353382 462218 388826 462454
rect 389062 462218 389146 462454
rect 389382 462218 424826 462454
rect 425062 462218 425146 462454
rect 425382 462218 460826 462454
rect 461062 462218 461146 462454
rect 461382 462218 496826 462454
rect 497062 462218 497146 462454
rect 497382 462218 532826 462454
rect 533062 462218 533146 462454
rect 533382 462218 568826 462454
rect 569062 462218 569146 462454
rect 569382 462218 591102 462454
rect 591338 462218 591422 462454
rect 591658 462218 592650 462454
rect -8726 462134 592650 462218
rect -8726 461898 -7734 462134
rect -7498 461898 -7414 462134
rect -7178 461898 28826 462134
rect 29062 461898 29146 462134
rect 29382 461898 64826 462134
rect 65062 461898 65146 462134
rect 65382 461898 100826 462134
rect 101062 461898 101146 462134
rect 101382 461898 136826 462134
rect 137062 461898 137146 462134
rect 137382 461898 172826 462134
rect 173062 461898 173146 462134
rect 173382 461898 208826 462134
rect 209062 461898 209146 462134
rect 209382 461898 244826 462134
rect 245062 461898 245146 462134
rect 245382 461898 280826 462134
rect 281062 461898 281146 462134
rect 281382 461898 316826 462134
rect 317062 461898 317146 462134
rect 317382 461898 352826 462134
rect 353062 461898 353146 462134
rect 353382 461898 388826 462134
rect 389062 461898 389146 462134
rect 389382 461898 424826 462134
rect 425062 461898 425146 462134
rect 425382 461898 460826 462134
rect 461062 461898 461146 462134
rect 461382 461898 496826 462134
rect 497062 461898 497146 462134
rect 497382 461898 532826 462134
rect 533062 461898 533146 462134
rect 533382 461898 568826 462134
rect 569062 461898 569146 462134
rect 569382 461898 591102 462134
rect 591338 461898 591422 462134
rect 591658 461898 592650 462134
rect -8726 461866 592650 461898
rect -8726 457954 592650 457986
rect -8726 457718 -6774 457954
rect -6538 457718 -6454 457954
rect -6218 457718 24326 457954
rect 24562 457718 24646 457954
rect 24882 457718 60326 457954
rect 60562 457718 60646 457954
rect 60882 457718 96326 457954
rect 96562 457718 96646 457954
rect 96882 457718 132326 457954
rect 132562 457718 132646 457954
rect 132882 457718 168326 457954
rect 168562 457718 168646 457954
rect 168882 457718 204326 457954
rect 204562 457718 204646 457954
rect 204882 457718 240326 457954
rect 240562 457718 240646 457954
rect 240882 457718 276326 457954
rect 276562 457718 276646 457954
rect 276882 457718 312326 457954
rect 312562 457718 312646 457954
rect 312882 457718 348326 457954
rect 348562 457718 348646 457954
rect 348882 457718 384326 457954
rect 384562 457718 384646 457954
rect 384882 457718 420326 457954
rect 420562 457718 420646 457954
rect 420882 457718 456326 457954
rect 456562 457718 456646 457954
rect 456882 457718 492326 457954
rect 492562 457718 492646 457954
rect 492882 457718 528326 457954
rect 528562 457718 528646 457954
rect 528882 457718 564326 457954
rect 564562 457718 564646 457954
rect 564882 457718 590142 457954
rect 590378 457718 590462 457954
rect 590698 457718 592650 457954
rect -8726 457634 592650 457718
rect -8726 457398 -6774 457634
rect -6538 457398 -6454 457634
rect -6218 457398 24326 457634
rect 24562 457398 24646 457634
rect 24882 457398 60326 457634
rect 60562 457398 60646 457634
rect 60882 457398 96326 457634
rect 96562 457398 96646 457634
rect 96882 457398 132326 457634
rect 132562 457398 132646 457634
rect 132882 457398 168326 457634
rect 168562 457398 168646 457634
rect 168882 457398 204326 457634
rect 204562 457398 204646 457634
rect 204882 457398 240326 457634
rect 240562 457398 240646 457634
rect 240882 457398 276326 457634
rect 276562 457398 276646 457634
rect 276882 457398 312326 457634
rect 312562 457398 312646 457634
rect 312882 457398 348326 457634
rect 348562 457398 348646 457634
rect 348882 457398 384326 457634
rect 384562 457398 384646 457634
rect 384882 457398 420326 457634
rect 420562 457398 420646 457634
rect 420882 457398 456326 457634
rect 456562 457398 456646 457634
rect 456882 457398 492326 457634
rect 492562 457398 492646 457634
rect 492882 457398 528326 457634
rect 528562 457398 528646 457634
rect 528882 457398 564326 457634
rect 564562 457398 564646 457634
rect 564882 457398 590142 457634
rect 590378 457398 590462 457634
rect 590698 457398 592650 457634
rect -8726 457366 592650 457398
rect -8726 453454 592650 453486
rect -8726 453218 -5814 453454
rect -5578 453218 -5494 453454
rect -5258 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 589182 453454
rect 589418 453218 589502 453454
rect 589738 453218 592650 453454
rect -8726 453134 592650 453218
rect -8726 452898 -5814 453134
rect -5578 452898 -5494 453134
rect -5258 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 589182 453134
rect 589418 452898 589502 453134
rect 589738 452898 592650 453134
rect -8726 452866 592650 452898
rect -8726 448954 592650 448986
rect -8726 448718 -4854 448954
rect -4618 448718 -4534 448954
rect -4298 448718 15326 448954
rect 15562 448718 15646 448954
rect 15882 448718 51326 448954
rect 51562 448718 51646 448954
rect 51882 448718 87326 448954
rect 87562 448718 87646 448954
rect 87882 448718 123326 448954
rect 123562 448718 123646 448954
rect 123882 448718 159326 448954
rect 159562 448718 159646 448954
rect 159882 448718 195326 448954
rect 195562 448718 195646 448954
rect 195882 448718 231326 448954
rect 231562 448718 231646 448954
rect 231882 448718 267326 448954
rect 267562 448718 267646 448954
rect 267882 448718 303326 448954
rect 303562 448718 303646 448954
rect 303882 448718 339326 448954
rect 339562 448718 339646 448954
rect 339882 448718 375326 448954
rect 375562 448718 375646 448954
rect 375882 448718 411326 448954
rect 411562 448718 411646 448954
rect 411882 448718 447326 448954
rect 447562 448718 447646 448954
rect 447882 448718 483326 448954
rect 483562 448718 483646 448954
rect 483882 448718 519326 448954
rect 519562 448718 519646 448954
rect 519882 448718 555326 448954
rect 555562 448718 555646 448954
rect 555882 448718 588222 448954
rect 588458 448718 588542 448954
rect 588778 448718 592650 448954
rect -8726 448634 592650 448718
rect -8726 448398 -4854 448634
rect -4618 448398 -4534 448634
rect -4298 448398 15326 448634
rect 15562 448398 15646 448634
rect 15882 448398 51326 448634
rect 51562 448398 51646 448634
rect 51882 448398 87326 448634
rect 87562 448398 87646 448634
rect 87882 448398 123326 448634
rect 123562 448398 123646 448634
rect 123882 448398 159326 448634
rect 159562 448398 159646 448634
rect 159882 448398 195326 448634
rect 195562 448398 195646 448634
rect 195882 448398 231326 448634
rect 231562 448398 231646 448634
rect 231882 448398 267326 448634
rect 267562 448398 267646 448634
rect 267882 448398 303326 448634
rect 303562 448398 303646 448634
rect 303882 448398 339326 448634
rect 339562 448398 339646 448634
rect 339882 448398 375326 448634
rect 375562 448398 375646 448634
rect 375882 448398 411326 448634
rect 411562 448398 411646 448634
rect 411882 448398 447326 448634
rect 447562 448398 447646 448634
rect 447882 448398 483326 448634
rect 483562 448398 483646 448634
rect 483882 448398 519326 448634
rect 519562 448398 519646 448634
rect 519882 448398 555326 448634
rect 555562 448398 555646 448634
rect 555882 448398 588222 448634
rect 588458 448398 588542 448634
rect 588778 448398 592650 448634
rect -8726 448366 592650 448398
rect -8726 444454 592650 444486
rect -8726 444218 -3894 444454
rect -3658 444218 -3574 444454
rect -3338 444218 10826 444454
rect 11062 444218 11146 444454
rect 11382 444218 46826 444454
rect 47062 444218 47146 444454
rect 47382 444218 82826 444454
rect 83062 444218 83146 444454
rect 83382 444218 118826 444454
rect 119062 444218 119146 444454
rect 119382 444218 154826 444454
rect 155062 444218 155146 444454
rect 155382 444218 190826 444454
rect 191062 444218 191146 444454
rect 191382 444218 226826 444454
rect 227062 444218 227146 444454
rect 227382 444218 262826 444454
rect 263062 444218 263146 444454
rect 263382 444218 298826 444454
rect 299062 444218 299146 444454
rect 299382 444218 334826 444454
rect 335062 444218 335146 444454
rect 335382 444218 370826 444454
rect 371062 444218 371146 444454
rect 371382 444218 406826 444454
rect 407062 444218 407146 444454
rect 407382 444218 442826 444454
rect 443062 444218 443146 444454
rect 443382 444218 478826 444454
rect 479062 444218 479146 444454
rect 479382 444218 514826 444454
rect 515062 444218 515146 444454
rect 515382 444218 550826 444454
rect 551062 444218 551146 444454
rect 551382 444218 587262 444454
rect 587498 444218 587582 444454
rect 587818 444218 592650 444454
rect -8726 444134 592650 444218
rect -8726 443898 -3894 444134
rect -3658 443898 -3574 444134
rect -3338 443898 10826 444134
rect 11062 443898 11146 444134
rect 11382 443898 46826 444134
rect 47062 443898 47146 444134
rect 47382 443898 82826 444134
rect 83062 443898 83146 444134
rect 83382 443898 118826 444134
rect 119062 443898 119146 444134
rect 119382 443898 154826 444134
rect 155062 443898 155146 444134
rect 155382 443898 190826 444134
rect 191062 443898 191146 444134
rect 191382 443898 226826 444134
rect 227062 443898 227146 444134
rect 227382 443898 262826 444134
rect 263062 443898 263146 444134
rect 263382 443898 298826 444134
rect 299062 443898 299146 444134
rect 299382 443898 334826 444134
rect 335062 443898 335146 444134
rect 335382 443898 370826 444134
rect 371062 443898 371146 444134
rect 371382 443898 406826 444134
rect 407062 443898 407146 444134
rect 407382 443898 442826 444134
rect 443062 443898 443146 444134
rect 443382 443898 478826 444134
rect 479062 443898 479146 444134
rect 479382 443898 514826 444134
rect 515062 443898 515146 444134
rect 515382 443898 550826 444134
rect 551062 443898 551146 444134
rect 551382 443898 587262 444134
rect 587498 443898 587582 444134
rect 587818 443898 592650 444134
rect -8726 443866 592650 443898
rect -8726 439954 592650 439986
rect -8726 439718 -2934 439954
rect -2698 439718 -2614 439954
rect -2378 439718 6326 439954
rect 6562 439718 6646 439954
rect 6882 439718 42326 439954
rect 42562 439718 42646 439954
rect 42882 439718 78326 439954
rect 78562 439718 78646 439954
rect 78882 439718 114326 439954
rect 114562 439718 114646 439954
rect 114882 439718 150326 439954
rect 150562 439718 150646 439954
rect 150882 439718 186326 439954
rect 186562 439718 186646 439954
rect 186882 439718 222326 439954
rect 222562 439718 222646 439954
rect 222882 439718 258326 439954
rect 258562 439718 258646 439954
rect 258882 439718 294326 439954
rect 294562 439718 294646 439954
rect 294882 439718 330326 439954
rect 330562 439718 330646 439954
rect 330882 439718 366326 439954
rect 366562 439718 366646 439954
rect 366882 439718 402326 439954
rect 402562 439718 402646 439954
rect 402882 439718 438326 439954
rect 438562 439718 438646 439954
rect 438882 439718 474326 439954
rect 474562 439718 474646 439954
rect 474882 439718 510326 439954
rect 510562 439718 510646 439954
rect 510882 439718 546326 439954
rect 546562 439718 546646 439954
rect 546882 439718 582326 439954
rect 582562 439718 582646 439954
rect 582882 439718 586302 439954
rect 586538 439718 586622 439954
rect 586858 439718 592650 439954
rect -8726 439634 592650 439718
rect -8726 439398 -2934 439634
rect -2698 439398 -2614 439634
rect -2378 439398 6326 439634
rect 6562 439398 6646 439634
rect 6882 439398 42326 439634
rect 42562 439398 42646 439634
rect 42882 439398 78326 439634
rect 78562 439398 78646 439634
rect 78882 439398 114326 439634
rect 114562 439398 114646 439634
rect 114882 439398 150326 439634
rect 150562 439398 150646 439634
rect 150882 439398 186326 439634
rect 186562 439398 186646 439634
rect 186882 439398 222326 439634
rect 222562 439398 222646 439634
rect 222882 439398 258326 439634
rect 258562 439398 258646 439634
rect 258882 439398 294326 439634
rect 294562 439398 294646 439634
rect 294882 439398 330326 439634
rect 330562 439398 330646 439634
rect 330882 439398 366326 439634
rect 366562 439398 366646 439634
rect 366882 439398 402326 439634
rect 402562 439398 402646 439634
rect 402882 439398 438326 439634
rect 438562 439398 438646 439634
rect 438882 439398 474326 439634
rect 474562 439398 474646 439634
rect 474882 439398 510326 439634
rect 510562 439398 510646 439634
rect 510882 439398 546326 439634
rect 546562 439398 546646 439634
rect 546882 439398 582326 439634
rect 582562 439398 582646 439634
rect 582882 439398 586302 439634
rect 586538 439398 586622 439634
rect 586858 439398 592650 439634
rect -8726 439366 592650 439398
rect -8726 435454 592650 435486
rect -8726 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 592650 435454
rect -8726 435134 592650 435218
rect -8726 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 592650 435134
rect -8726 434866 592650 434898
rect -8726 430954 592650 430986
rect -8726 430718 -8694 430954
rect -8458 430718 -8374 430954
rect -8138 430718 33326 430954
rect 33562 430718 33646 430954
rect 33882 430718 69326 430954
rect 69562 430718 69646 430954
rect 69882 430718 105326 430954
rect 105562 430718 105646 430954
rect 105882 430718 141326 430954
rect 141562 430718 141646 430954
rect 141882 430718 177326 430954
rect 177562 430718 177646 430954
rect 177882 430718 213326 430954
rect 213562 430718 213646 430954
rect 213882 430718 249326 430954
rect 249562 430718 249646 430954
rect 249882 430718 285326 430954
rect 285562 430718 285646 430954
rect 285882 430718 321326 430954
rect 321562 430718 321646 430954
rect 321882 430718 357326 430954
rect 357562 430718 357646 430954
rect 357882 430718 393326 430954
rect 393562 430718 393646 430954
rect 393882 430718 429326 430954
rect 429562 430718 429646 430954
rect 429882 430718 465326 430954
rect 465562 430718 465646 430954
rect 465882 430718 501326 430954
rect 501562 430718 501646 430954
rect 501882 430718 537326 430954
rect 537562 430718 537646 430954
rect 537882 430718 573326 430954
rect 573562 430718 573646 430954
rect 573882 430718 592062 430954
rect 592298 430718 592382 430954
rect 592618 430718 592650 430954
rect -8726 430634 592650 430718
rect -8726 430398 -8694 430634
rect -8458 430398 -8374 430634
rect -8138 430398 33326 430634
rect 33562 430398 33646 430634
rect 33882 430398 69326 430634
rect 69562 430398 69646 430634
rect 69882 430398 105326 430634
rect 105562 430398 105646 430634
rect 105882 430398 141326 430634
rect 141562 430398 141646 430634
rect 141882 430398 177326 430634
rect 177562 430398 177646 430634
rect 177882 430398 213326 430634
rect 213562 430398 213646 430634
rect 213882 430398 249326 430634
rect 249562 430398 249646 430634
rect 249882 430398 285326 430634
rect 285562 430398 285646 430634
rect 285882 430398 321326 430634
rect 321562 430398 321646 430634
rect 321882 430398 357326 430634
rect 357562 430398 357646 430634
rect 357882 430398 393326 430634
rect 393562 430398 393646 430634
rect 393882 430398 429326 430634
rect 429562 430398 429646 430634
rect 429882 430398 465326 430634
rect 465562 430398 465646 430634
rect 465882 430398 501326 430634
rect 501562 430398 501646 430634
rect 501882 430398 537326 430634
rect 537562 430398 537646 430634
rect 537882 430398 573326 430634
rect 573562 430398 573646 430634
rect 573882 430398 592062 430634
rect 592298 430398 592382 430634
rect 592618 430398 592650 430634
rect -8726 430366 592650 430398
rect -8726 426454 592650 426486
rect -8726 426218 -7734 426454
rect -7498 426218 -7414 426454
rect -7178 426218 28826 426454
rect 29062 426218 29146 426454
rect 29382 426218 64826 426454
rect 65062 426218 65146 426454
rect 65382 426218 100826 426454
rect 101062 426218 101146 426454
rect 101382 426218 136826 426454
rect 137062 426218 137146 426454
rect 137382 426218 172826 426454
rect 173062 426218 173146 426454
rect 173382 426218 208826 426454
rect 209062 426218 209146 426454
rect 209382 426218 244826 426454
rect 245062 426218 245146 426454
rect 245382 426218 280826 426454
rect 281062 426218 281146 426454
rect 281382 426218 316826 426454
rect 317062 426218 317146 426454
rect 317382 426218 352826 426454
rect 353062 426218 353146 426454
rect 353382 426218 388826 426454
rect 389062 426218 389146 426454
rect 389382 426218 424826 426454
rect 425062 426218 425146 426454
rect 425382 426218 460826 426454
rect 461062 426218 461146 426454
rect 461382 426218 496826 426454
rect 497062 426218 497146 426454
rect 497382 426218 532826 426454
rect 533062 426218 533146 426454
rect 533382 426218 568826 426454
rect 569062 426218 569146 426454
rect 569382 426218 591102 426454
rect 591338 426218 591422 426454
rect 591658 426218 592650 426454
rect -8726 426134 592650 426218
rect -8726 425898 -7734 426134
rect -7498 425898 -7414 426134
rect -7178 425898 28826 426134
rect 29062 425898 29146 426134
rect 29382 425898 64826 426134
rect 65062 425898 65146 426134
rect 65382 425898 100826 426134
rect 101062 425898 101146 426134
rect 101382 425898 136826 426134
rect 137062 425898 137146 426134
rect 137382 425898 172826 426134
rect 173062 425898 173146 426134
rect 173382 425898 208826 426134
rect 209062 425898 209146 426134
rect 209382 425898 244826 426134
rect 245062 425898 245146 426134
rect 245382 425898 280826 426134
rect 281062 425898 281146 426134
rect 281382 425898 316826 426134
rect 317062 425898 317146 426134
rect 317382 425898 352826 426134
rect 353062 425898 353146 426134
rect 353382 425898 388826 426134
rect 389062 425898 389146 426134
rect 389382 425898 424826 426134
rect 425062 425898 425146 426134
rect 425382 425898 460826 426134
rect 461062 425898 461146 426134
rect 461382 425898 496826 426134
rect 497062 425898 497146 426134
rect 497382 425898 532826 426134
rect 533062 425898 533146 426134
rect 533382 425898 568826 426134
rect 569062 425898 569146 426134
rect 569382 425898 591102 426134
rect 591338 425898 591422 426134
rect 591658 425898 592650 426134
rect -8726 425866 592650 425898
rect -8726 421954 592650 421986
rect -8726 421718 -6774 421954
rect -6538 421718 -6454 421954
rect -6218 421718 24326 421954
rect 24562 421718 24646 421954
rect 24882 421718 60326 421954
rect 60562 421718 60646 421954
rect 60882 421718 96326 421954
rect 96562 421718 96646 421954
rect 96882 421718 132326 421954
rect 132562 421718 132646 421954
rect 132882 421718 168326 421954
rect 168562 421718 168646 421954
rect 168882 421718 204326 421954
rect 204562 421718 204646 421954
rect 204882 421718 240326 421954
rect 240562 421718 240646 421954
rect 240882 421718 276326 421954
rect 276562 421718 276646 421954
rect 276882 421718 312326 421954
rect 312562 421718 312646 421954
rect 312882 421718 348326 421954
rect 348562 421718 348646 421954
rect 348882 421718 384326 421954
rect 384562 421718 384646 421954
rect 384882 421718 420326 421954
rect 420562 421718 420646 421954
rect 420882 421718 456326 421954
rect 456562 421718 456646 421954
rect 456882 421718 492326 421954
rect 492562 421718 492646 421954
rect 492882 421718 528326 421954
rect 528562 421718 528646 421954
rect 528882 421718 564326 421954
rect 564562 421718 564646 421954
rect 564882 421718 590142 421954
rect 590378 421718 590462 421954
rect 590698 421718 592650 421954
rect -8726 421634 592650 421718
rect -8726 421398 -6774 421634
rect -6538 421398 -6454 421634
rect -6218 421398 24326 421634
rect 24562 421398 24646 421634
rect 24882 421398 60326 421634
rect 60562 421398 60646 421634
rect 60882 421398 96326 421634
rect 96562 421398 96646 421634
rect 96882 421398 132326 421634
rect 132562 421398 132646 421634
rect 132882 421398 168326 421634
rect 168562 421398 168646 421634
rect 168882 421398 204326 421634
rect 204562 421398 204646 421634
rect 204882 421398 240326 421634
rect 240562 421398 240646 421634
rect 240882 421398 276326 421634
rect 276562 421398 276646 421634
rect 276882 421398 312326 421634
rect 312562 421398 312646 421634
rect 312882 421398 348326 421634
rect 348562 421398 348646 421634
rect 348882 421398 384326 421634
rect 384562 421398 384646 421634
rect 384882 421398 420326 421634
rect 420562 421398 420646 421634
rect 420882 421398 456326 421634
rect 456562 421398 456646 421634
rect 456882 421398 492326 421634
rect 492562 421398 492646 421634
rect 492882 421398 528326 421634
rect 528562 421398 528646 421634
rect 528882 421398 564326 421634
rect 564562 421398 564646 421634
rect 564882 421398 590142 421634
rect 590378 421398 590462 421634
rect 590698 421398 592650 421634
rect -8726 421366 592650 421398
rect -8726 417454 592650 417486
rect -8726 417218 -5814 417454
rect -5578 417218 -5494 417454
rect -5258 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 235826 417454
rect 236062 417218 236146 417454
rect 236382 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 343826 417454
rect 344062 417218 344146 417454
rect 344382 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 589182 417454
rect 589418 417218 589502 417454
rect 589738 417218 592650 417454
rect -8726 417134 592650 417218
rect -8726 416898 -5814 417134
rect -5578 416898 -5494 417134
rect -5258 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 235826 417134
rect 236062 416898 236146 417134
rect 236382 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 343826 417134
rect 344062 416898 344146 417134
rect 344382 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 589182 417134
rect 589418 416898 589502 417134
rect 589738 416898 592650 417134
rect -8726 416866 592650 416898
rect -8726 412954 592650 412986
rect -8726 412718 -4854 412954
rect -4618 412718 -4534 412954
rect -4298 412718 15326 412954
rect 15562 412718 15646 412954
rect 15882 412718 51326 412954
rect 51562 412718 51646 412954
rect 51882 412718 87326 412954
rect 87562 412718 87646 412954
rect 87882 412718 123326 412954
rect 123562 412718 123646 412954
rect 123882 412718 159326 412954
rect 159562 412718 159646 412954
rect 159882 412718 195326 412954
rect 195562 412718 195646 412954
rect 195882 412718 231326 412954
rect 231562 412718 231646 412954
rect 231882 412718 267326 412954
rect 267562 412718 267646 412954
rect 267882 412718 303326 412954
rect 303562 412718 303646 412954
rect 303882 412718 339326 412954
rect 339562 412718 339646 412954
rect 339882 412718 375326 412954
rect 375562 412718 375646 412954
rect 375882 412718 411326 412954
rect 411562 412718 411646 412954
rect 411882 412718 447326 412954
rect 447562 412718 447646 412954
rect 447882 412718 483326 412954
rect 483562 412718 483646 412954
rect 483882 412718 519326 412954
rect 519562 412718 519646 412954
rect 519882 412718 555326 412954
rect 555562 412718 555646 412954
rect 555882 412718 588222 412954
rect 588458 412718 588542 412954
rect 588778 412718 592650 412954
rect -8726 412634 592650 412718
rect -8726 412398 -4854 412634
rect -4618 412398 -4534 412634
rect -4298 412398 15326 412634
rect 15562 412398 15646 412634
rect 15882 412398 51326 412634
rect 51562 412398 51646 412634
rect 51882 412398 87326 412634
rect 87562 412398 87646 412634
rect 87882 412398 123326 412634
rect 123562 412398 123646 412634
rect 123882 412398 159326 412634
rect 159562 412398 159646 412634
rect 159882 412398 195326 412634
rect 195562 412398 195646 412634
rect 195882 412398 231326 412634
rect 231562 412398 231646 412634
rect 231882 412398 267326 412634
rect 267562 412398 267646 412634
rect 267882 412398 303326 412634
rect 303562 412398 303646 412634
rect 303882 412398 339326 412634
rect 339562 412398 339646 412634
rect 339882 412398 375326 412634
rect 375562 412398 375646 412634
rect 375882 412398 411326 412634
rect 411562 412398 411646 412634
rect 411882 412398 447326 412634
rect 447562 412398 447646 412634
rect 447882 412398 483326 412634
rect 483562 412398 483646 412634
rect 483882 412398 519326 412634
rect 519562 412398 519646 412634
rect 519882 412398 555326 412634
rect 555562 412398 555646 412634
rect 555882 412398 588222 412634
rect 588458 412398 588542 412634
rect 588778 412398 592650 412634
rect -8726 412366 592650 412398
rect -8726 408454 592650 408486
rect -8726 408218 -3894 408454
rect -3658 408218 -3574 408454
rect -3338 408218 10826 408454
rect 11062 408218 11146 408454
rect 11382 408218 46826 408454
rect 47062 408218 47146 408454
rect 47382 408218 82826 408454
rect 83062 408218 83146 408454
rect 83382 408218 118826 408454
rect 119062 408218 119146 408454
rect 119382 408218 154826 408454
rect 155062 408218 155146 408454
rect 155382 408218 190826 408454
rect 191062 408218 191146 408454
rect 191382 408218 226826 408454
rect 227062 408218 227146 408454
rect 227382 408218 262826 408454
rect 263062 408218 263146 408454
rect 263382 408218 298826 408454
rect 299062 408218 299146 408454
rect 299382 408218 334826 408454
rect 335062 408218 335146 408454
rect 335382 408218 370826 408454
rect 371062 408218 371146 408454
rect 371382 408218 406826 408454
rect 407062 408218 407146 408454
rect 407382 408218 442826 408454
rect 443062 408218 443146 408454
rect 443382 408218 478826 408454
rect 479062 408218 479146 408454
rect 479382 408218 514826 408454
rect 515062 408218 515146 408454
rect 515382 408218 550826 408454
rect 551062 408218 551146 408454
rect 551382 408218 587262 408454
rect 587498 408218 587582 408454
rect 587818 408218 592650 408454
rect -8726 408134 592650 408218
rect -8726 407898 -3894 408134
rect -3658 407898 -3574 408134
rect -3338 407898 10826 408134
rect 11062 407898 11146 408134
rect 11382 407898 46826 408134
rect 47062 407898 47146 408134
rect 47382 407898 82826 408134
rect 83062 407898 83146 408134
rect 83382 407898 118826 408134
rect 119062 407898 119146 408134
rect 119382 407898 154826 408134
rect 155062 407898 155146 408134
rect 155382 407898 190826 408134
rect 191062 407898 191146 408134
rect 191382 407898 226826 408134
rect 227062 407898 227146 408134
rect 227382 407898 262826 408134
rect 263062 407898 263146 408134
rect 263382 407898 298826 408134
rect 299062 407898 299146 408134
rect 299382 407898 334826 408134
rect 335062 407898 335146 408134
rect 335382 407898 370826 408134
rect 371062 407898 371146 408134
rect 371382 407898 406826 408134
rect 407062 407898 407146 408134
rect 407382 407898 442826 408134
rect 443062 407898 443146 408134
rect 443382 407898 478826 408134
rect 479062 407898 479146 408134
rect 479382 407898 514826 408134
rect 515062 407898 515146 408134
rect 515382 407898 550826 408134
rect 551062 407898 551146 408134
rect 551382 407898 587262 408134
rect 587498 407898 587582 408134
rect 587818 407898 592650 408134
rect -8726 407866 592650 407898
rect -8726 403954 592650 403986
rect -8726 403718 -2934 403954
rect -2698 403718 -2614 403954
rect -2378 403718 6326 403954
rect 6562 403718 6646 403954
rect 6882 403718 42326 403954
rect 42562 403718 42646 403954
rect 42882 403718 78326 403954
rect 78562 403718 78646 403954
rect 78882 403718 114326 403954
rect 114562 403718 114646 403954
rect 114882 403718 150326 403954
rect 150562 403718 150646 403954
rect 150882 403718 186326 403954
rect 186562 403718 186646 403954
rect 186882 403718 222326 403954
rect 222562 403718 222646 403954
rect 222882 403718 258326 403954
rect 258562 403718 258646 403954
rect 258882 403718 294326 403954
rect 294562 403718 294646 403954
rect 294882 403718 330326 403954
rect 330562 403718 330646 403954
rect 330882 403718 366326 403954
rect 366562 403718 366646 403954
rect 366882 403718 402326 403954
rect 402562 403718 402646 403954
rect 402882 403718 438326 403954
rect 438562 403718 438646 403954
rect 438882 403718 474326 403954
rect 474562 403718 474646 403954
rect 474882 403718 510326 403954
rect 510562 403718 510646 403954
rect 510882 403718 546326 403954
rect 546562 403718 546646 403954
rect 546882 403718 582326 403954
rect 582562 403718 582646 403954
rect 582882 403718 586302 403954
rect 586538 403718 586622 403954
rect 586858 403718 592650 403954
rect -8726 403634 592650 403718
rect -8726 403398 -2934 403634
rect -2698 403398 -2614 403634
rect -2378 403398 6326 403634
rect 6562 403398 6646 403634
rect 6882 403398 42326 403634
rect 42562 403398 42646 403634
rect 42882 403398 78326 403634
rect 78562 403398 78646 403634
rect 78882 403398 114326 403634
rect 114562 403398 114646 403634
rect 114882 403398 150326 403634
rect 150562 403398 150646 403634
rect 150882 403398 186326 403634
rect 186562 403398 186646 403634
rect 186882 403398 222326 403634
rect 222562 403398 222646 403634
rect 222882 403398 258326 403634
rect 258562 403398 258646 403634
rect 258882 403398 294326 403634
rect 294562 403398 294646 403634
rect 294882 403398 330326 403634
rect 330562 403398 330646 403634
rect 330882 403398 366326 403634
rect 366562 403398 366646 403634
rect 366882 403398 402326 403634
rect 402562 403398 402646 403634
rect 402882 403398 438326 403634
rect 438562 403398 438646 403634
rect 438882 403398 474326 403634
rect 474562 403398 474646 403634
rect 474882 403398 510326 403634
rect 510562 403398 510646 403634
rect 510882 403398 546326 403634
rect 546562 403398 546646 403634
rect 546882 403398 582326 403634
rect 582562 403398 582646 403634
rect 582882 403398 586302 403634
rect 586538 403398 586622 403634
rect 586858 403398 592650 403634
rect -8726 403366 592650 403398
rect -8726 399454 592650 399486
rect -8726 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 592650 399454
rect -8726 399134 592650 399218
rect -8726 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 592650 399134
rect -8726 398866 592650 398898
rect -8726 394954 592650 394986
rect -8726 394718 -8694 394954
rect -8458 394718 -8374 394954
rect -8138 394718 33326 394954
rect 33562 394718 33646 394954
rect 33882 394718 69326 394954
rect 69562 394718 69646 394954
rect 69882 394718 105326 394954
rect 105562 394718 105646 394954
rect 105882 394718 141326 394954
rect 141562 394718 141646 394954
rect 141882 394718 177326 394954
rect 177562 394718 177646 394954
rect 177882 394718 213326 394954
rect 213562 394718 213646 394954
rect 213882 394718 249326 394954
rect 249562 394718 249646 394954
rect 249882 394718 285326 394954
rect 285562 394718 285646 394954
rect 285882 394718 321326 394954
rect 321562 394718 321646 394954
rect 321882 394718 357326 394954
rect 357562 394718 357646 394954
rect 357882 394718 393326 394954
rect 393562 394718 393646 394954
rect 393882 394718 429326 394954
rect 429562 394718 429646 394954
rect 429882 394718 465326 394954
rect 465562 394718 465646 394954
rect 465882 394718 501326 394954
rect 501562 394718 501646 394954
rect 501882 394718 537326 394954
rect 537562 394718 537646 394954
rect 537882 394718 573326 394954
rect 573562 394718 573646 394954
rect 573882 394718 592062 394954
rect 592298 394718 592382 394954
rect 592618 394718 592650 394954
rect -8726 394634 592650 394718
rect -8726 394398 -8694 394634
rect -8458 394398 -8374 394634
rect -8138 394398 33326 394634
rect 33562 394398 33646 394634
rect 33882 394398 69326 394634
rect 69562 394398 69646 394634
rect 69882 394398 105326 394634
rect 105562 394398 105646 394634
rect 105882 394398 141326 394634
rect 141562 394398 141646 394634
rect 141882 394398 177326 394634
rect 177562 394398 177646 394634
rect 177882 394398 213326 394634
rect 213562 394398 213646 394634
rect 213882 394398 249326 394634
rect 249562 394398 249646 394634
rect 249882 394398 285326 394634
rect 285562 394398 285646 394634
rect 285882 394398 321326 394634
rect 321562 394398 321646 394634
rect 321882 394398 357326 394634
rect 357562 394398 357646 394634
rect 357882 394398 393326 394634
rect 393562 394398 393646 394634
rect 393882 394398 429326 394634
rect 429562 394398 429646 394634
rect 429882 394398 465326 394634
rect 465562 394398 465646 394634
rect 465882 394398 501326 394634
rect 501562 394398 501646 394634
rect 501882 394398 537326 394634
rect 537562 394398 537646 394634
rect 537882 394398 573326 394634
rect 573562 394398 573646 394634
rect 573882 394398 592062 394634
rect 592298 394398 592382 394634
rect 592618 394398 592650 394634
rect -8726 394366 592650 394398
rect -8726 390454 592650 390486
rect -8726 390218 -7734 390454
rect -7498 390218 -7414 390454
rect -7178 390218 28826 390454
rect 29062 390218 29146 390454
rect 29382 390218 64826 390454
rect 65062 390218 65146 390454
rect 65382 390218 100826 390454
rect 101062 390218 101146 390454
rect 101382 390218 136826 390454
rect 137062 390218 137146 390454
rect 137382 390218 172826 390454
rect 173062 390218 173146 390454
rect 173382 390218 208826 390454
rect 209062 390218 209146 390454
rect 209382 390218 244826 390454
rect 245062 390218 245146 390454
rect 245382 390218 280826 390454
rect 281062 390218 281146 390454
rect 281382 390218 316826 390454
rect 317062 390218 317146 390454
rect 317382 390218 352826 390454
rect 353062 390218 353146 390454
rect 353382 390218 388826 390454
rect 389062 390218 389146 390454
rect 389382 390218 424826 390454
rect 425062 390218 425146 390454
rect 425382 390218 460826 390454
rect 461062 390218 461146 390454
rect 461382 390218 496826 390454
rect 497062 390218 497146 390454
rect 497382 390218 532826 390454
rect 533062 390218 533146 390454
rect 533382 390218 568826 390454
rect 569062 390218 569146 390454
rect 569382 390218 591102 390454
rect 591338 390218 591422 390454
rect 591658 390218 592650 390454
rect -8726 390134 592650 390218
rect -8726 389898 -7734 390134
rect -7498 389898 -7414 390134
rect -7178 389898 28826 390134
rect 29062 389898 29146 390134
rect 29382 389898 64826 390134
rect 65062 389898 65146 390134
rect 65382 389898 100826 390134
rect 101062 389898 101146 390134
rect 101382 389898 136826 390134
rect 137062 389898 137146 390134
rect 137382 389898 172826 390134
rect 173062 389898 173146 390134
rect 173382 389898 208826 390134
rect 209062 389898 209146 390134
rect 209382 389898 244826 390134
rect 245062 389898 245146 390134
rect 245382 389898 280826 390134
rect 281062 389898 281146 390134
rect 281382 389898 316826 390134
rect 317062 389898 317146 390134
rect 317382 389898 352826 390134
rect 353062 389898 353146 390134
rect 353382 389898 388826 390134
rect 389062 389898 389146 390134
rect 389382 389898 424826 390134
rect 425062 389898 425146 390134
rect 425382 389898 460826 390134
rect 461062 389898 461146 390134
rect 461382 389898 496826 390134
rect 497062 389898 497146 390134
rect 497382 389898 532826 390134
rect 533062 389898 533146 390134
rect 533382 389898 568826 390134
rect 569062 389898 569146 390134
rect 569382 389898 591102 390134
rect 591338 389898 591422 390134
rect 591658 389898 592650 390134
rect -8726 389866 592650 389898
rect -8726 385954 592650 385986
rect -8726 385718 -6774 385954
rect -6538 385718 -6454 385954
rect -6218 385718 24326 385954
rect 24562 385718 24646 385954
rect 24882 385718 60326 385954
rect 60562 385718 60646 385954
rect 60882 385718 96326 385954
rect 96562 385718 96646 385954
rect 96882 385718 132326 385954
rect 132562 385718 132646 385954
rect 132882 385718 168326 385954
rect 168562 385718 168646 385954
rect 168882 385718 204326 385954
rect 204562 385718 204646 385954
rect 204882 385718 240326 385954
rect 240562 385718 240646 385954
rect 240882 385718 276326 385954
rect 276562 385718 276646 385954
rect 276882 385718 312326 385954
rect 312562 385718 312646 385954
rect 312882 385718 348326 385954
rect 348562 385718 348646 385954
rect 348882 385718 384326 385954
rect 384562 385718 384646 385954
rect 384882 385718 420326 385954
rect 420562 385718 420646 385954
rect 420882 385718 456326 385954
rect 456562 385718 456646 385954
rect 456882 385718 492326 385954
rect 492562 385718 492646 385954
rect 492882 385718 528326 385954
rect 528562 385718 528646 385954
rect 528882 385718 564326 385954
rect 564562 385718 564646 385954
rect 564882 385718 590142 385954
rect 590378 385718 590462 385954
rect 590698 385718 592650 385954
rect -8726 385634 592650 385718
rect -8726 385398 -6774 385634
rect -6538 385398 -6454 385634
rect -6218 385398 24326 385634
rect 24562 385398 24646 385634
rect 24882 385398 60326 385634
rect 60562 385398 60646 385634
rect 60882 385398 96326 385634
rect 96562 385398 96646 385634
rect 96882 385398 132326 385634
rect 132562 385398 132646 385634
rect 132882 385398 168326 385634
rect 168562 385398 168646 385634
rect 168882 385398 204326 385634
rect 204562 385398 204646 385634
rect 204882 385398 240326 385634
rect 240562 385398 240646 385634
rect 240882 385398 276326 385634
rect 276562 385398 276646 385634
rect 276882 385398 312326 385634
rect 312562 385398 312646 385634
rect 312882 385398 348326 385634
rect 348562 385398 348646 385634
rect 348882 385398 384326 385634
rect 384562 385398 384646 385634
rect 384882 385398 420326 385634
rect 420562 385398 420646 385634
rect 420882 385398 456326 385634
rect 456562 385398 456646 385634
rect 456882 385398 492326 385634
rect 492562 385398 492646 385634
rect 492882 385398 528326 385634
rect 528562 385398 528646 385634
rect 528882 385398 564326 385634
rect 564562 385398 564646 385634
rect 564882 385398 590142 385634
rect 590378 385398 590462 385634
rect 590698 385398 592650 385634
rect -8726 385366 592650 385398
rect -8726 381454 592650 381486
rect -8726 381218 -5814 381454
rect -5578 381218 -5494 381454
rect -5258 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 307826 381454
rect 308062 381218 308146 381454
rect 308382 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 589182 381454
rect 589418 381218 589502 381454
rect 589738 381218 592650 381454
rect -8726 381134 592650 381218
rect -8726 380898 -5814 381134
rect -5578 380898 -5494 381134
rect -5258 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 307826 381134
rect 308062 380898 308146 381134
rect 308382 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 589182 381134
rect 589418 380898 589502 381134
rect 589738 380898 592650 381134
rect -8726 380866 592650 380898
rect -8726 376954 592650 376986
rect -8726 376718 -4854 376954
rect -4618 376718 -4534 376954
rect -4298 376718 15326 376954
rect 15562 376718 15646 376954
rect 15882 376718 51326 376954
rect 51562 376718 51646 376954
rect 51882 376718 87326 376954
rect 87562 376718 87646 376954
rect 87882 376718 123326 376954
rect 123562 376718 123646 376954
rect 123882 376718 159326 376954
rect 159562 376718 159646 376954
rect 159882 376718 195326 376954
rect 195562 376718 195646 376954
rect 195882 376718 231326 376954
rect 231562 376718 231646 376954
rect 231882 376718 303326 376954
rect 303562 376718 303646 376954
rect 303882 376718 339326 376954
rect 339562 376718 339646 376954
rect 339882 376718 375326 376954
rect 375562 376718 375646 376954
rect 375882 376718 411326 376954
rect 411562 376718 411646 376954
rect 411882 376718 447326 376954
rect 447562 376718 447646 376954
rect 447882 376718 483326 376954
rect 483562 376718 483646 376954
rect 483882 376718 519326 376954
rect 519562 376718 519646 376954
rect 519882 376718 555326 376954
rect 555562 376718 555646 376954
rect 555882 376718 588222 376954
rect 588458 376718 588542 376954
rect 588778 376718 592650 376954
rect -8726 376634 592650 376718
rect -8726 376398 -4854 376634
rect -4618 376398 -4534 376634
rect -4298 376398 15326 376634
rect 15562 376398 15646 376634
rect 15882 376398 51326 376634
rect 51562 376398 51646 376634
rect 51882 376398 87326 376634
rect 87562 376398 87646 376634
rect 87882 376398 123326 376634
rect 123562 376398 123646 376634
rect 123882 376398 159326 376634
rect 159562 376398 159646 376634
rect 159882 376398 195326 376634
rect 195562 376398 195646 376634
rect 195882 376398 231326 376634
rect 231562 376398 231646 376634
rect 231882 376398 303326 376634
rect 303562 376398 303646 376634
rect 303882 376398 339326 376634
rect 339562 376398 339646 376634
rect 339882 376398 375326 376634
rect 375562 376398 375646 376634
rect 375882 376398 411326 376634
rect 411562 376398 411646 376634
rect 411882 376398 447326 376634
rect 447562 376398 447646 376634
rect 447882 376398 483326 376634
rect 483562 376398 483646 376634
rect 483882 376398 519326 376634
rect 519562 376398 519646 376634
rect 519882 376398 555326 376634
rect 555562 376398 555646 376634
rect 555882 376398 588222 376634
rect 588458 376398 588542 376634
rect 588778 376398 592650 376634
rect -8726 376366 592650 376398
rect -8726 372454 592650 372486
rect -8726 372218 -3894 372454
rect -3658 372218 -3574 372454
rect -3338 372218 10826 372454
rect 11062 372218 11146 372454
rect 11382 372218 46826 372454
rect 47062 372218 47146 372454
rect 47382 372218 82826 372454
rect 83062 372218 83146 372454
rect 83382 372218 118826 372454
rect 119062 372218 119146 372454
rect 119382 372218 154826 372454
rect 155062 372218 155146 372454
rect 155382 372218 190826 372454
rect 191062 372218 191146 372454
rect 191382 372218 226826 372454
rect 227062 372218 227146 372454
rect 227382 372218 334826 372454
rect 335062 372218 335146 372454
rect 335382 372218 370826 372454
rect 371062 372218 371146 372454
rect 371382 372218 406826 372454
rect 407062 372218 407146 372454
rect 407382 372218 442826 372454
rect 443062 372218 443146 372454
rect 443382 372218 478826 372454
rect 479062 372218 479146 372454
rect 479382 372218 514826 372454
rect 515062 372218 515146 372454
rect 515382 372218 550826 372454
rect 551062 372218 551146 372454
rect 551382 372218 587262 372454
rect 587498 372218 587582 372454
rect 587818 372218 592650 372454
rect -8726 372134 592650 372218
rect -8726 371898 -3894 372134
rect -3658 371898 -3574 372134
rect -3338 371898 10826 372134
rect 11062 371898 11146 372134
rect 11382 371898 46826 372134
rect 47062 371898 47146 372134
rect 47382 371898 82826 372134
rect 83062 371898 83146 372134
rect 83382 371898 118826 372134
rect 119062 371898 119146 372134
rect 119382 371898 154826 372134
rect 155062 371898 155146 372134
rect 155382 371898 190826 372134
rect 191062 371898 191146 372134
rect 191382 371898 226826 372134
rect 227062 371898 227146 372134
rect 227382 371898 334826 372134
rect 335062 371898 335146 372134
rect 335382 371898 370826 372134
rect 371062 371898 371146 372134
rect 371382 371898 406826 372134
rect 407062 371898 407146 372134
rect 407382 371898 442826 372134
rect 443062 371898 443146 372134
rect 443382 371898 478826 372134
rect 479062 371898 479146 372134
rect 479382 371898 514826 372134
rect 515062 371898 515146 372134
rect 515382 371898 550826 372134
rect 551062 371898 551146 372134
rect 551382 371898 587262 372134
rect 587498 371898 587582 372134
rect 587818 371898 592650 372134
rect -8726 371866 592650 371898
rect -8726 367954 592650 367986
rect -8726 367718 -2934 367954
rect -2698 367718 -2614 367954
rect -2378 367718 6326 367954
rect 6562 367718 6646 367954
rect 6882 367718 42326 367954
rect 42562 367718 42646 367954
rect 42882 367718 78326 367954
rect 78562 367718 78646 367954
rect 78882 367718 114326 367954
rect 114562 367718 114646 367954
rect 114882 367718 150326 367954
rect 150562 367718 150646 367954
rect 150882 367718 186326 367954
rect 186562 367718 186646 367954
rect 186882 367718 222326 367954
rect 222562 367718 222646 367954
rect 222882 367718 254610 367954
rect 254846 367718 285330 367954
rect 285566 367718 330326 367954
rect 330562 367718 330646 367954
rect 330882 367718 366326 367954
rect 366562 367718 366646 367954
rect 366882 367718 402326 367954
rect 402562 367718 402646 367954
rect 402882 367718 438326 367954
rect 438562 367718 438646 367954
rect 438882 367718 474326 367954
rect 474562 367718 474646 367954
rect 474882 367718 510326 367954
rect 510562 367718 510646 367954
rect 510882 367718 546326 367954
rect 546562 367718 546646 367954
rect 546882 367718 582326 367954
rect 582562 367718 582646 367954
rect 582882 367718 586302 367954
rect 586538 367718 586622 367954
rect 586858 367718 592650 367954
rect -8726 367634 592650 367718
rect -8726 367398 -2934 367634
rect -2698 367398 -2614 367634
rect -2378 367398 6326 367634
rect 6562 367398 6646 367634
rect 6882 367398 42326 367634
rect 42562 367398 42646 367634
rect 42882 367398 78326 367634
rect 78562 367398 78646 367634
rect 78882 367398 114326 367634
rect 114562 367398 114646 367634
rect 114882 367398 150326 367634
rect 150562 367398 150646 367634
rect 150882 367398 186326 367634
rect 186562 367398 186646 367634
rect 186882 367398 222326 367634
rect 222562 367398 222646 367634
rect 222882 367398 254610 367634
rect 254846 367398 285330 367634
rect 285566 367398 330326 367634
rect 330562 367398 330646 367634
rect 330882 367398 366326 367634
rect 366562 367398 366646 367634
rect 366882 367398 402326 367634
rect 402562 367398 402646 367634
rect 402882 367398 438326 367634
rect 438562 367398 438646 367634
rect 438882 367398 474326 367634
rect 474562 367398 474646 367634
rect 474882 367398 510326 367634
rect 510562 367398 510646 367634
rect 510882 367398 546326 367634
rect 546562 367398 546646 367634
rect 546882 367398 582326 367634
rect 582562 367398 582646 367634
rect 582882 367398 586302 367634
rect 586538 367398 586622 367634
rect 586858 367398 592650 367634
rect -8726 367366 592650 367398
rect -8726 363454 592650 363486
rect -8726 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 239250 363454
rect 239486 363218 269970 363454
rect 270206 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 592650 363454
rect -8726 363134 592650 363218
rect -8726 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 239250 363134
rect 239486 362898 269970 363134
rect 270206 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 592650 363134
rect -8726 362866 592650 362898
rect -8726 358954 592650 358986
rect -8726 358718 -8694 358954
rect -8458 358718 -8374 358954
rect -8138 358718 33326 358954
rect 33562 358718 33646 358954
rect 33882 358718 69326 358954
rect 69562 358718 69646 358954
rect 69882 358718 105326 358954
rect 105562 358718 105646 358954
rect 105882 358718 141326 358954
rect 141562 358718 141646 358954
rect 141882 358718 177326 358954
rect 177562 358718 177646 358954
rect 177882 358718 213326 358954
rect 213562 358718 213646 358954
rect 213882 358718 321326 358954
rect 321562 358718 321646 358954
rect 321882 358718 357326 358954
rect 357562 358718 357646 358954
rect 357882 358718 393326 358954
rect 393562 358718 393646 358954
rect 393882 358718 429326 358954
rect 429562 358718 429646 358954
rect 429882 358718 465326 358954
rect 465562 358718 465646 358954
rect 465882 358718 501326 358954
rect 501562 358718 501646 358954
rect 501882 358718 537326 358954
rect 537562 358718 537646 358954
rect 537882 358718 573326 358954
rect 573562 358718 573646 358954
rect 573882 358718 592062 358954
rect 592298 358718 592382 358954
rect 592618 358718 592650 358954
rect -8726 358634 592650 358718
rect -8726 358398 -8694 358634
rect -8458 358398 -8374 358634
rect -8138 358398 33326 358634
rect 33562 358398 33646 358634
rect 33882 358398 69326 358634
rect 69562 358398 69646 358634
rect 69882 358398 105326 358634
rect 105562 358398 105646 358634
rect 105882 358398 141326 358634
rect 141562 358398 141646 358634
rect 141882 358398 177326 358634
rect 177562 358398 177646 358634
rect 177882 358398 213326 358634
rect 213562 358398 213646 358634
rect 213882 358398 321326 358634
rect 321562 358398 321646 358634
rect 321882 358398 357326 358634
rect 357562 358398 357646 358634
rect 357882 358398 393326 358634
rect 393562 358398 393646 358634
rect 393882 358398 429326 358634
rect 429562 358398 429646 358634
rect 429882 358398 465326 358634
rect 465562 358398 465646 358634
rect 465882 358398 501326 358634
rect 501562 358398 501646 358634
rect 501882 358398 537326 358634
rect 537562 358398 537646 358634
rect 537882 358398 573326 358634
rect 573562 358398 573646 358634
rect 573882 358398 592062 358634
rect 592298 358398 592382 358634
rect 592618 358398 592650 358634
rect -8726 358366 592650 358398
rect -8726 354454 592650 354486
rect -8726 354218 -7734 354454
rect -7498 354218 -7414 354454
rect -7178 354218 28826 354454
rect 29062 354218 29146 354454
rect 29382 354218 64826 354454
rect 65062 354218 65146 354454
rect 65382 354218 100826 354454
rect 101062 354218 101146 354454
rect 101382 354218 136826 354454
rect 137062 354218 137146 354454
rect 137382 354218 172826 354454
rect 173062 354218 173146 354454
rect 173382 354218 208826 354454
rect 209062 354218 209146 354454
rect 209382 354218 316826 354454
rect 317062 354218 317146 354454
rect 317382 354218 352826 354454
rect 353062 354218 353146 354454
rect 353382 354218 388826 354454
rect 389062 354218 389146 354454
rect 389382 354218 424826 354454
rect 425062 354218 425146 354454
rect 425382 354218 460826 354454
rect 461062 354218 461146 354454
rect 461382 354218 496826 354454
rect 497062 354218 497146 354454
rect 497382 354218 532826 354454
rect 533062 354218 533146 354454
rect 533382 354218 568826 354454
rect 569062 354218 569146 354454
rect 569382 354218 591102 354454
rect 591338 354218 591422 354454
rect 591658 354218 592650 354454
rect -8726 354134 592650 354218
rect -8726 353898 -7734 354134
rect -7498 353898 -7414 354134
rect -7178 353898 28826 354134
rect 29062 353898 29146 354134
rect 29382 353898 64826 354134
rect 65062 353898 65146 354134
rect 65382 353898 100826 354134
rect 101062 353898 101146 354134
rect 101382 353898 136826 354134
rect 137062 353898 137146 354134
rect 137382 353898 172826 354134
rect 173062 353898 173146 354134
rect 173382 353898 208826 354134
rect 209062 353898 209146 354134
rect 209382 353898 316826 354134
rect 317062 353898 317146 354134
rect 317382 353898 352826 354134
rect 353062 353898 353146 354134
rect 353382 353898 388826 354134
rect 389062 353898 389146 354134
rect 389382 353898 424826 354134
rect 425062 353898 425146 354134
rect 425382 353898 460826 354134
rect 461062 353898 461146 354134
rect 461382 353898 496826 354134
rect 497062 353898 497146 354134
rect 497382 353898 532826 354134
rect 533062 353898 533146 354134
rect 533382 353898 568826 354134
rect 569062 353898 569146 354134
rect 569382 353898 591102 354134
rect 591338 353898 591422 354134
rect 591658 353898 592650 354134
rect -8726 353866 592650 353898
rect -8726 349954 592650 349986
rect -8726 349718 -6774 349954
rect -6538 349718 -6454 349954
rect -6218 349718 24326 349954
rect 24562 349718 24646 349954
rect 24882 349718 60326 349954
rect 60562 349718 60646 349954
rect 60882 349718 96326 349954
rect 96562 349718 96646 349954
rect 96882 349718 132326 349954
rect 132562 349718 132646 349954
rect 132882 349718 168326 349954
rect 168562 349718 168646 349954
rect 168882 349718 204326 349954
rect 204562 349718 204646 349954
rect 204882 349718 312326 349954
rect 312562 349718 312646 349954
rect 312882 349718 348326 349954
rect 348562 349718 348646 349954
rect 348882 349718 384326 349954
rect 384562 349718 384646 349954
rect 384882 349718 420326 349954
rect 420562 349718 420646 349954
rect 420882 349718 456326 349954
rect 456562 349718 456646 349954
rect 456882 349718 492326 349954
rect 492562 349718 492646 349954
rect 492882 349718 528326 349954
rect 528562 349718 528646 349954
rect 528882 349718 564326 349954
rect 564562 349718 564646 349954
rect 564882 349718 590142 349954
rect 590378 349718 590462 349954
rect 590698 349718 592650 349954
rect -8726 349634 592650 349718
rect -8726 349398 -6774 349634
rect -6538 349398 -6454 349634
rect -6218 349398 24326 349634
rect 24562 349398 24646 349634
rect 24882 349398 60326 349634
rect 60562 349398 60646 349634
rect 60882 349398 96326 349634
rect 96562 349398 96646 349634
rect 96882 349398 132326 349634
rect 132562 349398 132646 349634
rect 132882 349398 168326 349634
rect 168562 349398 168646 349634
rect 168882 349398 204326 349634
rect 204562 349398 204646 349634
rect 204882 349398 312326 349634
rect 312562 349398 312646 349634
rect 312882 349398 348326 349634
rect 348562 349398 348646 349634
rect 348882 349398 384326 349634
rect 384562 349398 384646 349634
rect 384882 349398 420326 349634
rect 420562 349398 420646 349634
rect 420882 349398 456326 349634
rect 456562 349398 456646 349634
rect 456882 349398 492326 349634
rect 492562 349398 492646 349634
rect 492882 349398 528326 349634
rect 528562 349398 528646 349634
rect 528882 349398 564326 349634
rect 564562 349398 564646 349634
rect 564882 349398 590142 349634
rect 590378 349398 590462 349634
rect 590698 349398 592650 349634
rect -8726 349366 592650 349398
rect -8726 345454 592650 345486
rect -8726 345218 -5814 345454
rect -5578 345218 -5494 345454
rect -5258 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 307826 345454
rect 308062 345218 308146 345454
rect 308382 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 589182 345454
rect 589418 345218 589502 345454
rect 589738 345218 592650 345454
rect -8726 345134 592650 345218
rect -8726 344898 -5814 345134
rect -5578 344898 -5494 345134
rect -5258 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 307826 345134
rect 308062 344898 308146 345134
rect 308382 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 589182 345134
rect 589418 344898 589502 345134
rect 589738 344898 592650 345134
rect -8726 344866 592650 344898
rect -8726 340954 592650 340986
rect -8726 340718 -4854 340954
rect -4618 340718 -4534 340954
rect -4298 340718 15326 340954
rect 15562 340718 15646 340954
rect 15882 340718 51326 340954
rect 51562 340718 51646 340954
rect 51882 340718 87326 340954
rect 87562 340718 87646 340954
rect 87882 340718 123326 340954
rect 123562 340718 123646 340954
rect 123882 340718 159326 340954
rect 159562 340718 159646 340954
rect 159882 340718 195326 340954
rect 195562 340718 195646 340954
rect 195882 340718 231326 340954
rect 231562 340718 231646 340954
rect 231882 340718 303326 340954
rect 303562 340718 303646 340954
rect 303882 340718 339326 340954
rect 339562 340718 339646 340954
rect 339882 340718 375326 340954
rect 375562 340718 375646 340954
rect 375882 340718 411326 340954
rect 411562 340718 411646 340954
rect 411882 340718 447326 340954
rect 447562 340718 447646 340954
rect 447882 340718 483326 340954
rect 483562 340718 483646 340954
rect 483882 340718 519326 340954
rect 519562 340718 519646 340954
rect 519882 340718 555326 340954
rect 555562 340718 555646 340954
rect 555882 340718 588222 340954
rect 588458 340718 588542 340954
rect 588778 340718 592650 340954
rect -8726 340634 592650 340718
rect -8726 340398 -4854 340634
rect -4618 340398 -4534 340634
rect -4298 340398 15326 340634
rect 15562 340398 15646 340634
rect 15882 340398 51326 340634
rect 51562 340398 51646 340634
rect 51882 340398 87326 340634
rect 87562 340398 87646 340634
rect 87882 340398 123326 340634
rect 123562 340398 123646 340634
rect 123882 340398 159326 340634
rect 159562 340398 159646 340634
rect 159882 340398 195326 340634
rect 195562 340398 195646 340634
rect 195882 340398 231326 340634
rect 231562 340398 231646 340634
rect 231882 340398 303326 340634
rect 303562 340398 303646 340634
rect 303882 340398 339326 340634
rect 339562 340398 339646 340634
rect 339882 340398 375326 340634
rect 375562 340398 375646 340634
rect 375882 340398 411326 340634
rect 411562 340398 411646 340634
rect 411882 340398 447326 340634
rect 447562 340398 447646 340634
rect 447882 340398 483326 340634
rect 483562 340398 483646 340634
rect 483882 340398 519326 340634
rect 519562 340398 519646 340634
rect 519882 340398 555326 340634
rect 555562 340398 555646 340634
rect 555882 340398 588222 340634
rect 588458 340398 588542 340634
rect 588778 340398 592650 340634
rect -8726 340366 592650 340398
rect -8726 336454 592650 336486
rect -8726 336218 -3894 336454
rect -3658 336218 -3574 336454
rect -3338 336218 10826 336454
rect 11062 336218 11146 336454
rect 11382 336218 46826 336454
rect 47062 336218 47146 336454
rect 47382 336218 82826 336454
rect 83062 336218 83146 336454
rect 83382 336218 118826 336454
rect 119062 336218 119146 336454
rect 119382 336218 154826 336454
rect 155062 336218 155146 336454
rect 155382 336218 190826 336454
rect 191062 336218 191146 336454
rect 191382 336218 226826 336454
rect 227062 336218 227146 336454
rect 227382 336218 334826 336454
rect 335062 336218 335146 336454
rect 335382 336218 370826 336454
rect 371062 336218 371146 336454
rect 371382 336218 406826 336454
rect 407062 336218 407146 336454
rect 407382 336218 442826 336454
rect 443062 336218 443146 336454
rect 443382 336218 478826 336454
rect 479062 336218 479146 336454
rect 479382 336218 514826 336454
rect 515062 336218 515146 336454
rect 515382 336218 550826 336454
rect 551062 336218 551146 336454
rect 551382 336218 587262 336454
rect 587498 336218 587582 336454
rect 587818 336218 592650 336454
rect -8726 336134 592650 336218
rect -8726 335898 -3894 336134
rect -3658 335898 -3574 336134
rect -3338 335898 10826 336134
rect 11062 335898 11146 336134
rect 11382 335898 46826 336134
rect 47062 335898 47146 336134
rect 47382 335898 82826 336134
rect 83062 335898 83146 336134
rect 83382 335898 118826 336134
rect 119062 335898 119146 336134
rect 119382 335898 154826 336134
rect 155062 335898 155146 336134
rect 155382 335898 190826 336134
rect 191062 335898 191146 336134
rect 191382 335898 226826 336134
rect 227062 335898 227146 336134
rect 227382 335898 334826 336134
rect 335062 335898 335146 336134
rect 335382 335898 370826 336134
rect 371062 335898 371146 336134
rect 371382 335898 406826 336134
rect 407062 335898 407146 336134
rect 407382 335898 442826 336134
rect 443062 335898 443146 336134
rect 443382 335898 478826 336134
rect 479062 335898 479146 336134
rect 479382 335898 514826 336134
rect 515062 335898 515146 336134
rect 515382 335898 550826 336134
rect 551062 335898 551146 336134
rect 551382 335898 587262 336134
rect 587498 335898 587582 336134
rect 587818 335898 592650 336134
rect -8726 335866 592650 335898
rect -8726 331954 592650 331986
rect -8726 331718 -2934 331954
rect -2698 331718 -2614 331954
rect -2378 331718 6326 331954
rect 6562 331718 6646 331954
rect 6882 331718 42326 331954
rect 42562 331718 42646 331954
rect 42882 331718 78326 331954
rect 78562 331718 78646 331954
rect 78882 331718 114326 331954
rect 114562 331718 114646 331954
rect 114882 331718 150326 331954
rect 150562 331718 150646 331954
rect 150882 331718 186326 331954
rect 186562 331718 186646 331954
rect 186882 331718 222326 331954
rect 222562 331718 222646 331954
rect 222882 331718 258326 331954
rect 258562 331718 258646 331954
rect 258882 331718 294326 331954
rect 294562 331718 294646 331954
rect 294882 331718 330326 331954
rect 330562 331718 330646 331954
rect 330882 331718 366326 331954
rect 366562 331718 366646 331954
rect 366882 331718 402326 331954
rect 402562 331718 402646 331954
rect 402882 331718 438326 331954
rect 438562 331718 438646 331954
rect 438882 331718 474326 331954
rect 474562 331718 474646 331954
rect 474882 331718 510326 331954
rect 510562 331718 510646 331954
rect 510882 331718 546326 331954
rect 546562 331718 546646 331954
rect 546882 331718 582326 331954
rect 582562 331718 582646 331954
rect 582882 331718 586302 331954
rect 586538 331718 586622 331954
rect 586858 331718 592650 331954
rect -8726 331634 592650 331718
rect -8726 331398 -2934 331634
rect -2698 331398 -2614 331634
rect -2378 331398 6326 331634
rect 6562 331398 6646 331634
rect 6882 331398 42326 331634
rect 42562 331398 42646 331634
rect 42882 331398 78326 331634
rect 78562 331398 78646 331634
rect 78882 331398 114326 331634
rect 114562 331398 114646 331634
rect 114882 331398 150326 331634
rect 150562 331398 150646 331634
rect 150882 331398 186326 331634
rect 186562 331398 186646 331634
rect 186882 331398 222326 331634
rect 222562 331398 222646 331634
rect 222882 331398 258326 331634
rect 258562 331398 258646 331634
rect 258882 331398 294326 331634
rect 294562 331398 294646 331634
rect 294882 331398 330326 331634
rect 330562 331398 330646 331634
rect 330882 331398 366326 331634
rect 366562 331398 366646 331634
rect 366882 331398 402326 331634
rect 402562 331398 402646 331634
rect 402882 331398 438326 331634
rect 438562 331398 438646 331634
rect 438882 331398 474326 331634
rect 474562 331398 474646 331634
rect 474882 331398 510326 331634
rect 510562 331398 510646 331634
rect 510882 331398 546326 331634
rect 546562 331398 546646 331634
rect 546882 331398 582326 331634
rect 582562 331398 582646 331634
rect 582882 331398 586302 331634
rect 586538 331398 586622 331634
rect 586858 331398 592650 331634
rect -8726 331366 592650 331398
rect -8726 327454 592650 327486
rect -8726 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 592650 327454
rect -8726 327134 592650 327218
rect -8726 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 592650 327134
rect -8726 326866 592650 326898
rect -8726 322954 592650 322986
rect -8726 322718 -8694 322954
rect -8458 322718 -8374 322954
rect -8138 322718 33326 322954
rect 33562 322718 33646 322954
rect 33882 322718 69326 322954
rect 69562 322718 69646 322954
rect 69882 322718 105326 322954
rect 105562 322718 105646 322954
rect 105882 322718 141326 322954
rect 141562 322718 141646 322954
rect 141882 322718 177326 322954
rect 177562 322718 177646 322954
rect 177882 322718 213326 322954
rect 213562 322718 213646 322954
rect 213882 322718 249326 322954
rect 249562 322718 249646 322954
rect 249882 322718 285326 322954
rect 285562 322718 285646 322954
rect 285882 322718 321326 322954
rect 321562 322718 321646 322954
rect 321882 322718 357326 322954
rect 357562 322718 357646 322954
rect 357882 322718 393326 322954
rect 393562 322718 393646 322954
rect 393882 322718 429326 322954
rect 429562 322718 429646 322954
rect 429882 322718 465326 322954
rect 465562 322718 465646 322954
rect 465882 322718 501326 322954
rect 501562 322718 501646 322954
rect 501882 322718 537326 322954
rect 537562 322718 537646 322954
rect 537882 322718 573326 322954
rect 573562 322718 573646 322954
rect 573882 322718 592062 322954
rect 592298 322718 592382 322954
rect 592618 322718 592650 322954
rect -8726 322634 592650 322718
rect -8726 322398 -8694 322634
rect -8458 322398 -8374 322634
rect -8138 322398 33326 322634
rect 33562 322398 33646 322634
rect 33882 322398 69326 322634
rect 69562 322398 69646 322634
rect 69882 322398 105326 322634
rect 105562 322398 105646 322634
rect 105882 322398 141326 322634
rect 141562 322398 141646 322634
rect 141882 322398 177326 322634
rect 177562 322398 177646 322634
rect 177882 322398 213326 322634
rect 213562 322398 213646 322634
rect 213882 322398 249326 322634
rect 249562 322398 249646 322634
rect 249882 322398 285326 322634
rect 285562 322398 285646 322634
rect 285882 322398 321326 322634
rect 321562 322398 321646 322634
rect 321882 322398 357326 322634
rect 357562 322398 357646 322634
rect 357882 322398 393326 322634
rect 393562 322398 393646 322634
rect 393882 322398 429326 322634
rect 429562 322398 429646 322634
rect 429882 322398 465326 322634
rect 465562 322398 465646 322634
rect 465882 322398 501326 322634
rect 501562 322398 501646 322634
rect 501882 322398 537326 322634
rect 537562 322398 537646 322634
rect 537882 322398 573326 322634
rect 573562 322398 573646 322634
rect 573882 322398 592062 322634
rect 592298 322398 592382 322634
rect 592618 322398 592650 322634
rect -8726 322366 592650 322398
rect -8726 318454 592650 318486
rect -8726 318218 -7734 318454
rect -7498 318218 -7414 318454
rect -7178 318218 28826 318454
rect 29062 318218 29146 318454
rect 29382 318218 64826 318454
rect 65062 318218 65146 318454
rect 65382 318218 100826 318454
rect 101062 318218 101146 318454
rect 101382 318218 136826 318454
rect 137062 318218 137146 318454
rect 137382 318218 172826 318454
rect 173062 318218 173146 318454
rect 173382 318218 208826 318454
rect 209062 318218 209146 318454
rect 209382 318218 244826 318454
rect 245062 318218 245146 318454
rect 245382 318218 280826 318454
rect 281062 318218 281146 318454
rect 281382 318218 316826 318454
rect 317062 318218 317146 318454
rect 317382 318218 352826 318454
rect 353062 318218 353146 318454
rect 353382 318218 388826 318454
rect 389062 318218 389146 318454
rect 389382 318218 424826 318454
rect 425062 318218 425146 318454
rect 425382 318218 460826 318454
rect 461062 318218 461146 318454
rect 461382 318218 496826 318454
rect 497062 318218 497146 318454
rect 497382 318218 532826 318454
rect 533062 318218 533146 318454
rect 533382 318218 568826 318454
rect 569062 318218 569146 318454
rect 569382 318218 591102 318454
rect 591338 318218 591422 318454
rect 591658 318218 592650 318454
rect -8726 318134 592650 318218
rect -8726 317898 -7734 318134
rect -7498 317898 -7414 318134
rect -7178 317898 28826 318134
rect 29062 317898 29146 318134
rect 29382 317898 64826 318134
rect 65062 317898 65146 318134
rect 65382 317898 100826 318134
rect 101062 317898 101146 318134
rect 101382 317898 136826 318134
rect 137062 317898 137146 318134
rect 137382 317898 172826 318134
rect 173062 317898 173146 318134
rect 173382 317898 208826 318134
rect 209062 317898 209146 318134
rect 209382 317898 244826 318134
rect 245062 317898 245146 318134
rect 245382 317898 280826 318134
rect 281062 317898 281146 318134
rect 281382 317898 316826 318134
rect 317062 317898 317146 318134
rect 317382 317898 352826 318134
rect 353062 317898 353146 318134
rect 353382 317898 388826 318134
rect 389062 317898 389146 318134
rect 389382 317898 424826 318134
rect 425062 317898 425146 318134
rect 425382 317898 460826 318134
rect 461062 317898 461146 318134
rect 461382 317898 496826 318134
rect 497062 317898 497146 318134
rect 497382 317898 532826 318134
rect 533062 317898 533146 318134
rect 533382 317898 568826 318134
rect 569062 317898 569146 318134
rect 569382 317898 591102 318134
rect 591338 317898 591422 318134
rect 591658 317898 592650 318134
rect -8726 317866 592650 317898
rect -8726 313954 592650 313986
rect -8726 313718 -6774 313954
rect -6538 313718 -6454 313954
rect -6218 313718 24326 313954
rect 24562 313718 24646 313954
rect 24882 313718 60326 313954
rect 60562 313718 60646 313954
rect 60882 313718 96326 313954
rect 96562 313718 96646 313954
rect 96882 313718 132326 313954
rect 132562 313718 132646 313954
rect 132882 313718 168326 313954
rect 168562 313718 168646 313954
rect 168882 313718 204326 313954
rect 204562 313718 204646 313954
rect 204882 313718 240326 313954
rect 240562 313718 240646 313954
rect 240882 313718 276326 313954
rect 276562 313718 276646 313954
rect 276882 313718 312326 313954
rect 312562 313718 312646 313954
rect 312882 313718 348326 313954
rect 348562 313718 348646 313954
rect 348882 313718 384326 313954
rect 384562 313718 384646 313954
rect 384882 313718 420326 313954
rect 420562 313718 420646 313954
rect 420882 313718 456326 313954
rect 456562 313718 456646 313954
rect 456882 313718 492326 313954
rect 492562 313718 492646 313954
rect 492882 313718 528326 313954
rect 528562 313718 528646 313954
rect 528882 313718 564326 313954
rect 564562 313718 564646 313954
rect 564882 313718 590142 313954
rect 590378 313718 590462 313954
rect 590698 313718 592650 313954
rect -8726 313634 592650 313718
rect -8726 313398 -6774 313634
rect -6538 313398 -6454 313634
rect -6218 313398 24326 313634
rect 24562 313398 24646 313634
rect 24882 313398 60326 313634
rect 60562 313398 60646 313634
rect 60882 313398 96326 313634
rect 96562 313398 96646 313634
rect 96882 313398 132326 313634
rect 132562 313398 132646 313634
rect 132882 313398 168326 313634
rect 168562 313398 168646 313634
rect 168882 313398 204326 313634
rect 204562 313398 204646 313634
rect 204882 313398 240326 313634
rect 240562 313398 240646 313634
rect 240882 313398 276326 313634
rect 276562 313398 276646 313634
rect 276882 313398 312326 313634
rect 312562 313398 312646 313634
rect 312882 313398 348326 313634
rect 348562 313398 348646 313634
rect 348882 313398 384326 313634
rect 384562 313398 384646 313634
rect 384882 313398 420326 313634
rect 420562 313398 420646 313634
rect 420882 313398 456326 313634
rect 456562 313398 456646 313634
rect 456882 313398 492326 313634
rect 492562 313398 492646 313634
rect 492882 313398 528326 313634
rect 528562 313398 528646 313634
rect 528882 313398 564326 313634
rect 564562 313398 564646 313634
rect 564882 313398 590142 313634
rect 590378 313398 590462 313634
rect 590698 313398 592650 313634
rect -8726 313366 592650 313398
rect -8726 309454 592650 309486
rect -8726 309218 -5814 309454
rect -5578 309218 -5494 309454
rect -5258 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 235826 309454
rect 236062 309218 236146 309454
rect 236382 309218 271826 309454
rect 272062 309218 272146 309454
rect 272382 309218 307826 309454
rect 308062 309218 308146 309454
rect 308382 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 589182 309454
rect 589418 309218 589502 309454
rect 589738 309218 592650 309454
rect -8726 309134 592650 309218
rect -8726 308898 -5814 309134
rect -5578 308898 -5494 309134
rect -5258 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 235826 309134
rect 236062 308898 236146 309134
rect 236382 308898 271826 309134
rect 272062 308898 272146 309134
rect 272382 308898 307826 309134
rect 308062 308898 308146 309134
rect 308382 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 589182 309134
rect 589418 308898 589502 309134
rect 589738 308898 592650 309134
rect -8726 308866 592650 308898
rect -8726 304954 592650 304986
rect -8726 304718 -4854 304954
rect -4618 304718 -4534 304954
rect -4298 304718 15326 304954
rect 15562 304718 15646 304954
rect 15882 304718 51326 304954
rect 51562 304718 51646 304954
rect 51882 304718 87326 304954
rect 87562 304718 87646 304954
rect 87882 304718 123326 304954
rect 123562 304718 123646 304954
rect 123882 304718 159326 304954
rect 159562 304718 159646 304954
rect 159882 304718 195326 304954
rect 195562 304718 195646 304954
rect 195882 304718 231326 304954
rect 231562 304718 231646 304954
rect 231882 304718 267326 304954
rect 267562 304718 267646 304954
rect 267882 304718 303326 304954
rect 303562 304718 303646 304954
rect 303882 304718 339326 304954
rect 339562 304718 339646 304954
rect 339882 304718 375326 304954
rect 375562 304718 375646 304954
rect 375882 304718 411326 304954
rect 411562 304718 411646 304954
rect 411882 304718 447326 304954
rect 447562 304718 447646 304954
rect 447882 304718 483326 304954
rect 483562 304718 483646 304954
rect 483882 304718 519326 304954
rect 519562 304718 519646 304954
rect 519882 304718 555326 304954
rect 555562 304718 555646 304954
rect 555882 304718 588222 304954
rect 588458 304718 588542 304954
rect 588778 304718 592650 304954
rect -8726 304634 592650 304718
rect -8726 304398 -4854 304634
rect -4618 304398 -4534 304634
rect -4298 304398 15326 304634
rect 15562 304398 15646 304634
rect 15882 304398 51326 304634
rect 51562 304398 51646 304634
rect 51882 304398 87326 304634
rect 87562 304398 87646 304634
rect 87882 304398 123326 304634
rect 123562 304398 123646 304634
rect 123882 304398 159326 304634
rect 159562 304398 159646 304634
rect 159882 304398 195326 304634
rect 195562 304398 195646 304634
rect 195882 304398 231326 304634
rect 231562 304398 231646 304634
rect 231882 304398 267326 304634
rect 267562 304398 267646 304634
rect 267882 304398 303326 304634
rect 303562 304398 303646 304634
rect 303882 304398 339326 304634
rect 339562 304398 339646 304634
rect 339882 304398 375326 304634
rect 375562 304398 375646 304634
rect 375882 304398 411326 304634
rect 411562 304398 411646 304634
rect 411882 304398 447326 304634
rect 447562 304398 447646 304634
rect 447882 304398 483326 304634
rect 483562 304398 483646 304634
rect 483882 304398 519326 304634
rect 519562 304398 519646 304634
rect 519882 304398 555326 304634
rect 555562 304398 555646 304634
rect 555882 304398 588222 304634
rect 588458 304398 588542 304634
rect 588778 304398 592650 304634
rect -8726 304366 592650 304398
rect -8726 300454 592650 300486
rect -8726 300218 -3894 300454
rect -3658 300218 -3574 300454
rect -3338 300218 10826 300454
rect 11062 300218 11146 300454
rect 11382 300218 46826 300454
rect 47062 300218 47146 300454
rect 47382 300218 82826 300454
rect 83062 300218 83146 300454
rect 83382 300218 118826 300454
rect 119062 300218 119146 300454
rect 119382 300218 154826 300454
rect 155062 300218 155146 300454
rect 155382 300218 190826 300454
rect 191062 300218 191146 300454
rect 191382 300218 226826 300454
rect 227062 300218 227146 300454
rect 227382 300218 262826 300454
rect 263062 300218 263146 300454
rect 263382 300218 298826 300454
rect 299062 300218 299146 300454
rect 299382 300218 334826 300454
rect 335062 300218 335146 300454
rect 335382 300218 370826 300454
rect 371062 300218 371146 300454
rect 371382 300218 406826 300454
rect 407062 300218 407146 300454
rect 407382 300218 442826 300454
rect 443062 300218 443146 300454
rect 443382 300218 478826 300454
rect 479062 300218 479146 300454
rect 479382 300218 514826 300454
rect 515062 300218 515146 300454
rect 515382 300218 550826 300454
rect 551062 300218 551146 300454
rect 551382 300218 587262 300454
rect 587498 300218 587582 300454
rect 587818 300218 592650 300454
rect -8726 300134 592650 300218
rect -8726 299898 -3894 300134
rect -3658 299898 -3574 300134
rect -3338 299898 10826 300134
rect 11062 299898 11146 300134
rect 11382 299898 46826 300134
rect 47062 299898 47146 300134
rect 47382 299898 82826 300134
rect 83062 299898 83146 300134
rect 83382 299898 118826 300134
rect 119062 299898 119146 300134
rect 119382 299898 154826 300134
rect 155062 299898 155146 300134
rect 155382 299898 190826 300134
rect 191062 299898 191146 300134
rect 191382 299898 226826 300134
rect 227062 299898 227146 300134
rect 227382 299898 262826 300134
rect 263062 299898 263146 300134
rect 263382 299898 298826 300134
rect 299062 299898 299146 300134
rect 299382 299898 334826 300134
rect 335062 299898 335146 300134
rect 335382 299898 370826 300134
rect 371062 299898 371146 300134
rect 371382 299898 406826 300134
rect 407062 299898 407146 300134
rect 407382 299898 442826 300134
rect 443062 299898 443146 300134
rect 443382 299898 478826 300134
rect 479062 299898 479146 300134
rect 479382 299898 514826 300134
rect 515062 299898 515146 300134
rect 515382 299898 550826 300134
rect 551062 299898 551146 300134
rect 551382 299898 587262 300134
rect 587498 299898 587582 300134
rect 587818 299898 592650 300134
rect -8726 299866 592650 299898
rect -8726 295954 592650 295986
rect -8726 295718 -2934 295954
rect -2698 295718 -2614 295954
rect -2378 295718 6326 295954
rect 6562 295718 6646 295954
rect 6882 295718 42326 295954
rect 42562 295718 42646 295954
rect 42882 295718 78326 295954
rect 78562 295718 78646 295954
rect 78882 295718 114326 295954
rect 114562 295718 114646 295954
rect 114882 295718 150326 295954
rect 150562 295718 150646 295954
rect 150882 295718 186326 295954
rect 186562 295718 186646 295954
rect 186882 295718 222326 295954
rect 222562 295718 222646 295954
rect 222882 295718 258326 295954
rect 258562 295718 258646 295954
rect 258882 295718 294326 295954
rect 294562 295718 294646 295954
rect 294882 295718 330326 295954
rect 330562 295718 330646 295954
rect 330882 295718 366326 295954
rect 366562 295718 366646 295954
rect 366882 295718 402326 295954
rect 402562 295718 402646 295954
rect 402882 295718 438326 295954
rect 438562 295718 438646 295954
rect 438882 295718 474326 295954
rect 474562 295718 474646 295954
rect 474882 295718 510326 295954
rect 510562 295718 510646 295954
rect 510882 295718 546326 295954
rect 546562 295718 546646 295954
rect 546882 295718 582326 295954
rect 582562 295718 582646 295954
rect 582882 295718 586302 295954
rect 586538 295718 586622 295954
rect 586858 295718 592650 295954
rect -8726 295634 592650 295718
rect -8726 295398 -2934 295634
rect -2698 295398 -2614 295634
rect -2378 295398 6326 295634
rect 6562 295398 6646 295634
rect 6882 295398 42326 295634
rect 42562 295398 42646 295634
rect 42882 295398 78326 295634
rect 78562 295398 78646 295634
rect 78882 295398 114326 295634
rect 114562 295398 114646 295634
rect 114882 295398 150326 295634
rect 150562 295398 150646 295634
rect 150882 295398 186326 295634
rect 186562 295398 186646 295634
rect 186882 295398 222326 295634
rect 222562 295398 222646 295634
rect 222882 295398 258326 295634
rect 258562 295398 258646 295634
rect 258882 295398 294326 295634
rect 294562 295398 294646 295634
rect 294882 295398 330326 295634
rect 330562 295398 330646 295634
rect 330882 295398 366326 295634
rect 366562 295398 366646 295634
rect 366882 295398 402326 295634
rect 402562 295398 402646 295634
rect 402882 295398 438326 295634
rect 438562 295398 438646 295634
rect 438882 295398 474326 295634
rect 474562 295398 474646 295634
rect 474882 295398 510326 295634
rect 510562 295398 510646 295634
rect 510882 295398 546326 295634
rect 546562 295398 546646 295634
rect 546882 295398 582326 295634
rect 582562 295398 582646 295634
rect 582882 295398 586302 295634
rect 586538 295398 586622 295634
rect 586858 295398 592650 295634
rect -8726 295366 592650 295398
rect -8726 291454 592650 291486
rect -8726 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 592650 291454
rect -8726 291134 592650 291218
rect -8726 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 592650 291134
rect -8726 290866 592650 290898
rect -8726 286954 592650 286986
rect -8726 286718 -8694 286954
rect -8458 286718 -8374 286954
rect -8138 286718 33326 286954
rect 33562 286718 33646 286954
rect 33882 286718 69326 286954
rect 69562 286718 69646 286954
rect 69882 286718 105326 286954
rect 105562 286718 105646 286954
rect 105882 286718 141326 286954
rect 141562 286718 141646 286954
rect 141882 286718 177326 286954
rect 177562 286718 177646 286954
rect 177882 286718 213326 286954
rect 213562 286718 213646 286954
rect 213882 286718 249326 286954
rect 249562 286718 249646 286954
rect 249882 286718 285326 286954
rect 285562 286718 285646 286954
rect 285882 286718 321326 286954
rect 321562 286718 321646 286954
rect 321882 286718 357326 286954
rect 357562 286718 357646 286954
rect 357882 286718 393326 286954
rect 393562 286718 393646 286954
rect 393882 286718 429326 286954
rect 429562 286718 429646 286954
rect 429882 286718 465326 286954
rect 465562 286718 465646 286954
rect 465882 286718 501326 286954
rect 501562 286718 501646 286954
rect 501882 286718 537326 286954
rect 537562 286718 537646 286954
rect 537882 286718 573326 286954
rect 573562 286718 573646 286954
rect 573882 286718 592062 286954
rect 592298 286718 592382 286954
rect 592618 286718 592650 286954
rect -8726 286634 592650 286718
rect -8726 286398 -8694 286634
rect -8458 286398 -8374 286634
rect -8138 286398 33326 286634
rect 33562 286398 33646 286634
rect 33882 286398 69326 286634
rect 69562 286398 69646 286634
rect 69882 286398 105326 286634
rect 105562 286398 105646 286634
rect 105882 286398 141326 286634
rect 141562 286398 141646 286634
rect 141882 286398 177326 286634
rect 177562 286398 177646 286634
rect 177882 286398 213326 286634
rect 213562 286398 213646 286634
rect 213882 286398 249326 286634
rect 249562 286398 249646 286634
rect 249882 286398 285326 286634
rect 285562 286398 285646 286634
rect 285882 286398 321326 286634
rect 321562 286398 321646 286634
rect 321882 286398 357326 286634
rect 357562 286398 357646 286634
rect 357882 286398 393326 286634
rect 393562 286398 393646 286634
rect 393882 286398 429326 286634
rect 429562 286398 429646 286634
rect 429882 286398 465326 286634
rect 465562 286398 465646 286634
rect 465882 286398 501326 286634
rect 501562 286398 501646 286634
rect 501882 286398 537326 286634
rect 537562 286398 537646 286634
rect 537882 286398 573326 286634
rect 573562 286398 573646 286634
rect 573882 286398 592062 286634
rect 592298 286398 592382 286634
rect 592618 286398 592650 286634
rect -8726 286366 592650 286398
rect -8726 282454 592650 282486
rect -8726 282218 -7734 282454
rect -7498 282218 -7414 282454
rect -7178 282218 28826 282454
rect 29062 282218 29146 282454
rect 29382 282218 64826 282454
rect 65062 282218 65146 282454
rect 65382 282218 100826 282454
rect 101062 282218 101146 282454
rect 101382 282218 136826 282454
rect 137062 282218 137146 282454
rect 137382 282218 172826 282454
rect 173062 282218 173146 282454
rect 173382 282218 208826 282454
rect 209062 282218 209146 282454
rect 209382 282218 244826 282454
rect 245062 282218 245146 282454
rect 245382 282218 280826 282454
rect 281062 282218 281146 282454
rect 281382 282218 316826 282454
rect 317062 282218 317146 282454
rect 317382 282218 352826 282454
rect 353062 282218 353146 282454
rect 353382 282218 388826 282454
rect 389062 282218 389146 282454
rect 389382 282218 424826 282454
rect 425062 282218 425146 282454
rect 425382 282218 460826 282454
rect 461062 282218 461146 282454
rect 461382 282218 496826 282454
rect 497062 282218 497146 282454
rect 497382 282218 532826 282454
rect 533062 282218 533146 282454
rect 533382 282218 568826 282454
rect 569062 282218 569146 282454
rect 569382 282218 591102 282454
rect 591338 282218 591422 282454
rect 591658 282218 592650 282454
rect -8726 282134 592650 282218
rect -8726 281898 -7734 282134
rect -7498 281898 -7414 282134
rect -7178 281898 28826 282134
rect 29062 281898 29146 282134
rect 29382 281898 64826 282134
rect 65062 281898 65146 282134
rect 65382 281898 100826 282134
rect 101062 281898 101146 282134
rect 101382 281898 136826 282134
rect 137062 281898 137146 282134
rect 137382 281898 172826 282134
rect 173062 281898 173146 282134
rect 173382 281898 208826 282134
rect 209062 281898 209146 282134
rect 209382 281898 244826 282134
rect 245062 281898 245146 282134
rect 245382 281898 280826 282134
rect 281062 281898 281146 282134
rect 281382 281898 316826 282134
rect 317062 281898 317146 282134
rect 317382 281898 352826 282134
rect 353062 281898 353146 282134
rect 353382 281898 388826 282134
rect 389062 281898 389146 282134
rect 389382 281898 424826 282134
rect 425062 281898 425146 282134
rect 425382 281898 460826 282134
rect 461062 281898 461146 282134
rect 461382 281898 496826 282134
rect 497062 281898 497146 282134
rect 497382 281898 532826 282134
rect 533062 281898 533146 282134
rect 533382 281898 568826 282134
rect 569062 281898 569146 282134
rect 569382 281898 591102 282134
rect 591338 281898 591422 282134
rect 591658 281898 592650 282134
rect -8726 281866 592650 281898
rect -8726 277954 592650 277986
rect -8726 277718 -6774 277954
rect -6538 277718 -6454 277954
rect -6218 277718 24326 277954
rect 24562 277718 24646 277954
rect 24882 277718 60326 277954
rect 60562 277718 60646 277954
rect 60882 277718 96326 277954
rect 96562 277718 96646 277954
rect 96882 277718 132326 277954
rect 132562 277718 132646 277954
rect 132882 277718 168326 277954
rect 168562 277718 168646 277954
rect 168882 277718 204326 277954
rect 204562 277718 204646 277954
rect 204882 277718 240326 277954
rect 240562 277718 240646 277954
rect 240882 277718 276326 277954
rect 276562 277718 276646 277954
rect 276882 277718 312326 277954
rect 312562 277718 312646 277954
rect 312882 277718 348326 277954
rect 348562 277718 348646 277954
rect 348882 277718 384326 277954
rect 384562 277718 384646 277954
rect 384882 277718 420326 277954
rect 420562 277718 420646 277954
rect 420882 277718 456326 277954
rect 456562 277718 456646 277954
rect 456882 277718 492326 277954
rect 492562 277718 492646 277954
rect 492882 277718 528326 277954
rect 528562 277718 528646 277954
rect 528882 277718 564326 277954
rect 564562 277718 564646 277954
rect 564882 277718 590142 277954
rect 590378 277718 590462 277954
rect 590698 277718 592650 277954
rect -8726 277634 592650 277718
rect -8726 277398 -6774 277634
rect -6538 277398 -6454 277634
rect -6218 277398 24326 277634
rect 24562 277398 24646 277634
rect 24882 277398 60326 277634
rect 60562 277398 60646 277634
rect 60882 277398 96326 277634
rect 96562 277398 96646 277634
rect 96882 277398 132326 277634
rect 132562 277398 132646 277634
rect 132882 277398 168326 277634
rect 168562 277398 168646 277634
rect 168882 277398 204326 277634
rect 204562 277398 204646 277634
rect 204882 277398 240326 277634
rect 240562 277398 240646 277634
rect 240882 277398 276326 277634
rect 276562 277398 276646 277634
rect 276882 277398 312326 277634
rect 312562 277398 312646 277634
rect 312882 277398 348326 277634
rect 348562 277398 348646 277634
rect 348882 277398 384326 277634
rect 384562 277398 384646 277634
rect 384882 277398 420326 277634
rect 420562 277398 420646 277634
rect 420882 277398 456326 277634
rect 456562 277398 456646 277634
rect 456882 277398 492326 277634
rect 492562 277398 492646 277634
rect 492882 277398 528326 277634
rect 528562 277398 528646 277634
rect 528882 277398 564326 277634
rect 564562 277398 564646 277634
rect 564882 277398 590142 277634
rect 590378 277398 590462 277634
rect 590698 277398 592650 277634
rect -8726 277366 592650 277398
rect -8726 273454 592650 273486
rect -8726 273218 -5814 273454
rect -5578 273218 -5494 273454
rect -5258 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 91826 273454
rect 92062 273218 92146 273454
rect 92382 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 199826 273454
rect 200062 273218 200146 273454
rect 200382 273218 235826 273454
rect 236062 273218 236146 273454
rect 236382 273218 271826 273454
rect 272062 273218 272146 273454
rect 272382 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 589182 273454
rect 589418 273218 589502 273454
rect 589738 273218 592650 273454
rect -8726 273134 592650 273218
rect -8726 272898 -5814 273134
rect -5578 272898 -5494 273134
rect -5258 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 91826 273134
rect 92062 272898 92146 273134
rect 92382 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 199826 273134
rect 200062 272898 200146 273134
rect 200382 272898 235826 273134
rect 236062 272898 236146 273134
rect 236382 272898 271826 273134
rect 272062 272898 272146 273134
rect 272382 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 589182 273134
rect 589418 272898 589502 273134
rect 589738 272898 592650 273134
rect -8726 272866 592650 272898
rect -8726 268954 592650 268986
rect -8726 268718 -4854 268954
rect -4618 268718 -4534 268954
rect -4298 268718 15326 268954
rect 15562 268718 15646 268954
rect 15882 268718 51326 268954
rect 51562 268718 51646 268954
rect 51882 268718 87326 268954
rect 87562 268718 87646 268954
rect 87882 268718 123326 268954
rect 123562 268718 123646 268954
rect 123882 268718 159326 268954
rect 159562 268718 159646 268954
rect 159882 268718 195326 268954
rect 195562 268718 195646 268954
rect 195882 268718 231326 268954
rect 231562 268718 231646 268954
rect 231882 268718 267326 268954
rect 267562 268718 267646 268954
rect 267882 268718 303326 268954
rect 303562 268718 303646 268954
rect 303882 268718 339326 268954
rect 339562 268718 339646 268954
rect 339882 268718 375326 268954
rect 375562 268718 375646 268954
rect 375882 268718 411326 268954
rect 411562 268718 411646 268954
rect 411882 268718 447326 268954
rect 447562 268718 447646 268954
rect 447882 268718 483326 268954
rect 483562 268718 483646 268954
rect 483882 268718 519326 268954
rect 519562 268718 519646 268954
rect 519882 268718 555326 268954
rect 555562 268718 555646 268954
rect 555882 268718 588222 268954
rect 588458 268718 588542 268954
rect 588778 268718 592650 268954
rect -8726 268634 592650 268718
rect -8726 268398 -4854 268634
rect -4618 268398 -4534 268634
rect -4298 268398 15326 268634
rect 15562 268398 15646 268634
rect 15882 268398 51326 268634
rect 51562 268398 51646 268634
rect 51882 268398 87326 268634
rect 87562 268398 87646 268634
rect 87882 268398 123326 268634
rect 123562 268398 123646 268634
rect 123882 268398 159326 268634
rect 159562 268398 159646 268634
rect 159882 268398 195326 268634
rect 195562 268398 195646 268634
rect 195882 268398 231326 268634
rect 231562 268398 231646 268634
rect 231882 268398 267326 268634
rect 267562 268398 267646 268634
rect 267882 268398 303326 268634
rect 303562 268398 303646 268634
rect 303882 268398 339326 268634
rect 339562 268398 339646 268634
rect 339882 268398 375326 268634
rect 375562 268398 375646 268634
rect 375882 268398 411326 268634
rect 411562 268398 411646 268634
rect 411882 268398 447326 268634
rect 447562 268398 447646 268634
rect 447882 268398 483326 268634
rect 483562 268398 483646 268634
rect 483882 268398 519326 268634
rect 519562 268398 519646 268634
rect 519882 268398 555326 268634
rect 555562 268398 555646 268634
rect 555882 268398 588222 268634
rect 588458 268398 588542 268634
rect 588778 268398 592650 268634
rect -8726 268366 592650 268398
rect -8726 264454 592650 264486
rect -8726 264218 -3894 264454
rect -3658 264218 -3574 264454
rect -3338 264218 10826 264454
rect 11062 264218 11146 264454
rect 11382 264218 46826 264454
rect 47062 264218 47146 264454
rect 47382 264218 82826 264454
rect 83062 264218 83146 264454
rect 83382 264218 118826 264454
rect 119062 264218 119146 264454
rect 119382 264218 154826 264454
rect 155062 264218 155146 264454
rect 155382 264218 190826 264454
rect 191062 264218 191146 264454
rect 191382 264218 226826 264454
rect 227062 264218 227146 264454
rect 227382 264218 262826 264454
rect 263062 264218 263146 264454
rect 263382 264218 298826 264454
rect 299062 264218 299146 264454
rect 299382 264218 334826 264454
rect 335062 264218 335146 264454
rect 335382 264218 370826 264454
rect 371062 264218 371146 264454
rect 371382 264218 406826 264454
rect 407062 264218 407146 264454
rect 407382 264218 442826 264454
rect 443062 264218 443146 264454
rect 443382 264218 478826 264454
rect 479062 264218 479146 264454
rect 479382 264218 514826 264454
rect 515062 264218 515146 264454
rect 515382 264218 550826 264454
rect 551062 264218 551146 264454
rect 551382 264218 587262 264454
rect 587498 264218 587582 264454
rect 587818 264218 592650 264454
rect -8726 264134 592650 264218
rect -8726 263898 -3894 264134
rect -3658 263898 -3574 264134
rect -3338 263898 10826 264134
rect 11062 263898 11146 264134
rect 11382 263898 46826 264134
rect 47062 263898 47146 264134
rect 47382 263898 82826 264134
rect 83062 263898 83146 264134
rect 83382 263898 118826 264134
rect 119062 263898 119146 264134
rect 119382 263898 154826 264134
rect 155062 263898 155146 264134
rect 155382 263898 190826 264134
rect 191062 263898 191146 264134
rect 191382 263898 226826 264134
rect 227062 263898 227146 264134
rect 227382 263898 262826 264134
rect 263062 263898 263146 264134
rect 263382 263898 298826 264134
rect 299062 263898 299146 264134
rect 299382 263898 334826 264134
rect 335062 263898 335146 264134
rect 335382 263898 370826 264134
rect 371062 263898 371146 264134
rect 371382 263898 406826 264134
rect 407062 263898 407146 264134
rect 407382 263898 442826 264134
rect 443062 263898 443146 264134
rect 443382 263898 478826 264134
rect 479062 263898 479146 264134
rect 479382 263898 514826 264134
rect 515062 263898 515146 264134
rect 515382 263898 550826 264134
rect 551062 263898 551146 264134
rect 551382 263898 587262 264134
rect 587498 263898 587582 264134
rect 587818 263898 592650 264134
rect -8726 263866 592650 263898
rect -8726 259954 592650 259986
rect -8726 259718 -2934 259954
rect -2698 259718 -2614 259954
rect -2378 259718 6326 259954
rect 6562 259718 6646 259954
rect 6882 259718 42326 259954
rect 42562 259718 42646 259954
rect 42882 259718 78326 259954
rect 78562 259718 78646 259954
rect 78882 259718 114326 259954
rect 114562 259718 114646 259954
rect 114882 259718 150326 259954
rect 150562 259718 150646 259954
rect 150882 259718 186326 259954
rect 186562 259718 186646 259954
rect 186882 259718 222326 259954
rect 222562 259718 222646 259954
rect 222882 259718 258326 259954
rect 258562 259718 258646 259954
rect 258882 259718 294326 259954
rect 294562 259718 294646 259954
rect 294882 259718 330326 259954
rect 330562 259718 330646 259954
rect 330882 259718 366326 259954
rect 366562 259718 366646 259954
rect 366882 259718 402326 259954
rect 402562 259718 402646 259954
rect 402882 259718 438326 259954
rect 438562 259718 438646 259954
rect 438882 259718 474326 259954
rect 474562 259718 474646 259954
rect 474882 259718 510326 259954
rect 510562 259718 510646 259954
rect 510882 259718 546326 259954
rect 546562 259718 546646 259954
rect 546882 259718 582326 259954
rect 582562 259718 582646 259954
rect 582882 259718 586302 259954
rect 586538 259718 586622 259954
rect 586858 259718 592650 259954
rect -8726 259634 592650 259718
rect -8726 259398 -2934 259634
rect -2698 259398 -2614 259634
rect -2378 259398 6326 259634
rect 6562 259398 6646 259634
rect 6882 259398 42326 259634
rect 42562 259398 42646 259634
rect 42882 259398 78326 259634
rect 78562 259398 78646 259634
rect 78882 259398 114326 259634
rect 114562 259398 114646 259634
rect 114882 259398 150326 259634
rect 150562 259398 150646 259634
rect 150882 259398 186326 259634
rect 186562 259398 186646 259634
rect 186882 259398 222326 259634
rect 222562 259398 222646 259634
rect 222882 259398 258326 259634
rect 258562 259398 258646 259634
rect 258882 259398 294326 259634
rect 294562 259398 294646 259634
rect 294882 259398 330326 259634
rect 330562 259398 330646 259634
rect 330882 259398 366326 259634
rect 366562 259398 366646 259634
rect 366882 259398 402326 259634
rect 402562 259398 402646 259634
rect 402882 259398 438326 259634
rect 438562 259398 438646 259634
rect 438882 259398 474326 259634
rect 474562 259398 474646 259634
rect 474882 259398 510326 259634
rect 510562 259398 510646 259634
rect 510882 259398 546326 259634
rect 546562 259398 546646 259634
rect 546882 259398 582326 259634
rect 582562 259398 582646 259634
rect 582882 259398 586302 259634
rect 586538 259398 586622 259634
rect 586858 259398 592650 259634
rect -8726 259366 592650 259398
rect -8726 255454 592650 255486
rect -8726 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 592650 255454
rect -8726 255134 592650 255218
rect -8726 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 592650 255134
rect -8726 254866 592650 254898
rect -8726 250954 592650 250986
rect -8726 250718 -8694 250954
rect -8458 250718 -8374 250954
rect -8138 250718 33326 250954
rect 33562 250718 33646 250954
rect 33882 250718 69326 250954
rect 69562 250718 69646 250954
rect 69882 250718 105326 250954
rect 105562 250718 105646 250954
rect 105882 250718 141326 250954
rect 141562 250718 141646 250954
rect 141882 250718 177326 250954
rect 177562 250718 177646 250954
rect 177882 250718 213326 250954
rect 213562 250718 213646 250954
rect 213882 250718 249326 250954
rect 249562 250718 249646 250954
rect 249882 250718 285326 250954
rect 285562 250718 285646 250954
rect 285882 250718 321326 250954
rect 321562 250718 321646 250954
rect 321882 250718 357326 250954
rect 357562 250718 357646 250954
rect 357882 250718 393326 250954
rect 393562 250718 393646 250954
rect 393882 250718 429326 250954
rect 429562 250718 429646 250954
rect 429882 250718 465326 250954
rect 465562 250718 465646 250954
rect 465882 250718 501326 250954
rect 501562 250718 501646 250954
rect 501882 250718 537326 250954
rect 537562 250718 537646 250954
rect 537882 250718 573326 250954
rect 573562 250718 573646 250954
rect 573882 250718 592062 250954
rect 592298 250718 592382 250954
rect 592618 250718 592650 250954
rect -8726 250634 592650 250718
rect -8726 250398 -8694 250634
rect -8458 250398 -8374 250634
rect -8138 250398 33326 250634
rect 33562 250398 33646 250634
rect 33882 250398 69326 250634
rect 69562 250398 69646 250634
rect 69882 250398 105326 250634
rect 105562 250398 105646 250634
rect 105882 250398 141326 250634
rect 141562 250398 141646 250634
rect 141882 250398 177326 250634
rect 177562 250398 177646 250634
rect 177882 250398 213326 250634
rect 213562 250398 213646 250634
rect 213882 250398 249326 250634
rect 249562 250398 249646 250634
rect 249882 250398 285326 250634
rect 285562 250398 285646 250634
rect 285882 250398 321326 250634
rect 321562 250398 321646 250634
rect 321882 250398 357326 250634
rect 357562 250398 357646 250634
rect 357882 250398 393326 250634
rect 393562 250398 393646 250634
rect 393882 250398 429326 250634
rect 429562 250398 429646 250634
rect 429882 250398 465326 250634
rect 465562 250398 465646 250634
rect 465882 250398 501326 250634
rect 501562 250398 501646 250634
rect 501882 250398 537326 250634
rect 537562 250398 537646 250634
rect 537882 250398 573326 250634
rect 573562 250398 573646 250634
rect 573882 250398 592062 250634
rect 592298 250398 592382 250634
rect 592618 250398 592650 250634
rect -8726 250366 592650 250398
rect -8726 246454 592650 246486
rect -8726 246218 -7734 246454
rect -7498 246218 -7414 246454
rect -7178 246218 28826 246454
rect 29062 246218 29146 246454
rect 29382 246218 64826 246454
rect 65062 246218 65146 246454
rect 65382 246218 100826 246454
rect 101062 246218 101146 246454
rect 101382 246218 136826 246454
rect 137062 246218 137146 246454
rect 137382 246218 172826 246454
rect 173062 246218 173146 246454
rect 173382 246218 208826 246454
rect 209062 246218 209146 246454
rect 209382 246218 244826 246454
rect 245062 246218 245146 246454
rect 245382 246218 280826 246454
rect 281062 246218 281146 246454
rect 281382 246218 316826 246454
rect 317062 246218 317146 246454
rect 317382 246218 352826 246454
rect 353062 246218 353146 246454
rect 353382 246218 388826 246454
rect 389062 246218 389146 246454
rect 389382 246218 424826 246454
rect 425062 246218 425146 246454
rect 425382 246218 460826 246454
rect 461062 246218 461146 246454
rect 461382 246218 496826 246454
rect 497062 246218 497146 246454
rect 497382 246218 532826 246454
rect 533062 246218 533146 246454
rect 533382 246218 568826 246454
rect 569062 246218 569146 246454
rect 569382 246218 591102 246454
rect 591338 246218 591422 246454
rect 591658 246218 592650 246454
rect -8726 246134 592650 246218
rect -8726 245898 -7734 246134
rect -7498 245898 -7414 246134
rect -7178 245898 28826 246134
rect 29062 245898 29146 246134
rect 29382 245898 64826 246134
rect 65062 245898 65146 246134
rect 65382 245898 100826 246134
rect 101062 245898 101146 246134
rect 101382 245898 136826 246134
rect 137062 245898 137146 246134
rect 137382 245898 172826 246134
rect 173062 245898 173146 246134
rect 173382 245898 208826 246134
rect 209062 245898 209146 246134
rect 209382 245898 244826 246134
rect 245062 245898 245146 246134
rect 245382 245898 280826 246134
rect 281062 245898 281146 246134
rect 281382 245898 316826 246134
rect 317062 245898 317146 246134
rect 317382 245898 352826 246134
rect 353062 245898 353146 246134
rect 353382 245898 388826 246134
rect 389062 245898 389146 246134
rect 389382 245898 424826 246134
rect 425062 245898 425146 246134
rect 425382 245898 460826 246134
rect 461062 245898 461146 246134
rect 461382 245898 496826 246134
rect 497062 245898 497146 246134
rect 497382 245898 532826 246134
rect 533062 245898 533146 246134
rect 533382 245898 568826 246134
rect 569062 245898 569146 246134
rect 569382 245898 591102 246134
rect 591338 245898 591422 246134
rect 591658 245898 592650 246134
rect -8726 245866 592650 245898
rect -8726 241954 592650 241986
rect -8726 241718 -6774 241954
rect -6538 241718 -6454 241954
rect -6218 241718 24326 241954
rect 24562 241718 24646 241954
rect 24882 241718 60326 241954
rect 60562 241718 60646 241954
rect 60882 241718 96326 241954
rect 96562 241718 96646 241954
rect 96882 241718 132326 241954
rect 132562 241718 132646 241954
rect 132882 241718 168326 241954
rect 168562 241718 168646 241954
rect 168882 241718 204326 241954
rect 204562 241718 204646 241954
rect 204882 241718 240326 241954
rect 240562 241718 240646 241954
rect 240882 241718 276326 241954
rect 276562 241718 276646 241954
rect 276882 241718 312326 241954
rect 312562 241718 312646 241954
rect 312882 241718 348326 241954
rect 348562 241718 348646 241954
rect 348882 241718 384326 241954
rect 384562 241718 384646 241954
rect 384882 241718 420326 241954
rect 420562 241718 420646 241954
rect 420882 241718 456326 241954
rect 456562 241718 456646 241954
rect 456882 241718 492326 241954
rect 492562 241718 492646 241954
rect 492882 241718 528326 241954
rect 528562 241718 528646 241954
rect 528882 241718 564326 241954
rect 564562 241718 564646 241954
rect 564882 241718 590142 241954
rect 590378 241718 590462 241954
rect 590698 241718 592650 241954
rect -8726 241634 592650 241718
rect -8726 241398 -6774 241634
rect -6538 241398 -6454 241634
rect -6218 241398 24326 241634
rect 24562 241398 24646 241634
rect 24882 241398 60326 241634
rect 60562 241398 60646 241634
rect 60882 241398 96326 241634
rect 96562 241398 96646 241634
rect 96882 241398 132326 241634
rect 132562 241398 132646 241634
rect 132882 241398 168326 241634
rect 168562 241398 168646 241634
rect 168882 241398 204326 241634
rect 204562 241398 204646 241634
rect 204882 241398 240326 241634
rect 240562 241398 240646 241634
rect 240882 241398 276326 241634
rect 276562 241398 276646 241634
rect 276882 241398 312326 241634
rect 312562 241398 312646 241634
rect 312882 241398 348326 241634
rect 348562 241398 348646 241634
rect 348882 241398 384326 241634
rect 384562 241398 384646 241634
rect 384882 241398 420326 241634
rect 420562 241398 420646 241634
rect 420882 241398 456326 241634
rect 456562 241398 456646 241634
rect 456882 241398 492326 241634
rect 492562 241398 492646 241634
rect 492882 241398 528326 241634
rect 528562 241398 528646 241634
rect 528882 241398 564326 241634
rect 564562 241398 564646 241634
rect 564882 241398 590142 241634
rect 590378 241398 590462 241634
rect 590698 241398 592650 241634
rect -8726 241366 592650 241398
rect -8726 237454 592650 237486
rect -8726 237218 -5814 237454
rect -5578 237218 -5494 237454
rect -5258 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 127826 237454
rect 128062 237218 128146 237454
rect 128382 237218 163826 237454
rect 164062 237218 164146 237454
rect 164382 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 235826 237454
rect 236062 237218 236146 237454
rect 236382 237218 271826 237454
rect 272062 237218 272146 237454
rect 272382 237218 307826 237454
rect 308062 237218 308146 237454
rect 308382 237218 343826 237454
rect 344062 237218 344146 237454
rect 344382 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 589182 237454
rect 589418 237218 589502 237454
rect 589738 237218 592650 237454
rect -8726 237134 592650 237218
rect -8726 236898 -5814 237134
rect -5578 236898 -5494 237134
rect -5258 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 127826 237134
rect 128062 236898 128146 237134
rect 128382 236898 163826 237134
rect 164062 236898 164146 237134
rect 164382 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 235826 237134
rect 236062 236898 236146 237134
rect 236382 236898 271826 237134
rect 272062 236898 272146 237134
rect 272382 236898 307826 237134
rect 308062 236898 308146 237134
rect 308382 236898 343826 237134
rect 344062 236898 344146 237134
rect 344382 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 589182 237134
rect 589418 236898 589502 237134
rect 589738 236898 592650 237134
rect -8726 236866 592650 236898
rect -8726 232954 592650 232986
rect -8726 232718 -4854 232954
rect -4618 232718 -4534 232954
rect -4298 232718 15326 232954
rect 15562 232718 15646 232954
rect 15882 232718 51326 232954
rect 51562 232718 51646 232954
rect 51882 232718 87326 232954
rect 87562 232718 87646 232954
rect 87882 232718 123326 232954
rect 123562 232718 123646 232954
rect 123882 232718 159326 232954
rect 159562 232718 159646 232954
rect 159882 232718 195326 232954
rect 195562 232718 195646 232954
rect 195882 232718 231326 232954
rect 231562 232718 231646 232954
rect 231882 232718 267326 232954
rect 267562 232718 267646 232954
rect 267882 232718 303326 232954
rect 303562 232718 303646 232954
rect 303882 232718 339326 232954
rect 339562 232718 339646 232954
rect 339882 232718 375326 232954
rect 375562 232718 375646 232954
rect 375882 232718 411326 232954
rect 411562 232718 411646 232954
rect 411882 232718 447326 232954
rect 447562 232718 447646 232954
rect 447882 232718 483326 232954
rect 483562 232718 483646 232954
rect 483882 232718 519326 232954
rect 519562 232718 519646 232954
rect 519882 232718 555326 232954
rect 555562 232718 555646 232954
rect 555882 232718 588222 232954
rect 588458 232718 588542 232954
rect 588778 232718 592650 232954
rect -8726 232634 592650 232718
rect -8726 232398 -4854 232634
rect -4618 232398 -4534 232634
rect -4298 232398 15326 232634
rect 15562 232398 15646 232634
rect 15882 232398 51326 232634
rect 51562 232398 51646 232634
rect 51882 232398 87326 232634
rect 87562 232398 87646 232634
rect 87882 232398 123326 232634
rect 123562 232398 123646 232634
rect 123882 232398 159326 232634
rect 159562 232398 159646 232634
rect 159882 232398 195326 232634
rect 195562 232398 195646 232634
rect 195882 232398 231326 232634
rect 231562 232398 231646 232634
rect 231882 232398 267326 232634
rect 267562 232398 267646 232634
rect 267882 232398 303326 232634
rect 303562 232398 303646 232634
rect 303882 232398 339326 232634
rect 339562 232398 339646 232634
rect 339882 232398 375326 232634
rect 375562 232398 375646 232634
rect 375882 232398 411326 232634
rect 411562 232398 411646 232634
rect 411882 232398 447326 232634
rect 447562 232398 447646 232634
rect 447882 232398 483326 232634
rect 483562 232398 483646 232634
rect 483882 232398 519326 232634
rect 519562 232398 519646 232634
rect 519882 232398 555326 232634
rect 555562 232398 555646 232634
rect 555882 232398 588222 232634
rect 588458 232398 588542 232634
rect 588778 232398 592650 232634
rect -8726 232366 592650 232398
rect -8726 228454 592650 228486
rect -8726 228218 -3894 228454
rect -3658 228218 -3574 228454
rect -3338 228218 10826 228454
rect 11062 228218 11146 228454
rect 11382 228218 46826 228454
rect 47062 228218 47146 228454
rect 47382 228218 82826 228454
rect 83062 228218 83146 228454
rect 83382 228218 118826 228454
rect 119062 228218 119146 228454
rect 119382 228218 154826 228454
rect 155062 228218 155146 228454
rect 155382 228218 190826 228454
rect 191062 228218 191146 228454
rect 191382 228218 226826 228454
rect 227062 228218 227146 228454
rect 227382 228218 262826 228454
rect 263062 228218 263146 228454
rect 263382 228218 298826 228454
rect 299062 228218 299146 228454
rect 299382 228218 334826 228454
rect 335062 228218 335146 228454
rect 335382 228218 370826 228454
rect 371062 228218 371146 228454
rect 371382 228218 406826 228454
rect 407062 228218 407146 228454
rect 407382 228218 442826 228454
rect 443062 228218 443146 228454
rect 443382 228218 478826 228454
rect 479062 228218 479146 228454
rect 479382 228218 514826 228454
rect 515062 228218 515146 228454
rect 515382 228218 550826 228454
rect 551062 228218 551146 228454
rect 551382 228218 587262 228454
rect 587498 228218 587582 228454
rect 587818 228218 592650 228454
rect -8726 228134 592650 228218
rect -8726 227898 -3894 228134
rect -3658 227898 -3574 228134
rect -3338 227898 10826 228134
rect 11062 227898 11146 228134
rect 11382 227898 46826 228134
rect 47062 227898 47146 228134
rect 47382 227898 82826 228134
rect 83062 227898 83146 228134
rect 83382 227898 118826 228134
rect 119062 227898 119146 228134
rect 119382 227898 154826 228134
rect 155062 227898 155146 228134
rect 155382 227898 190826 228134
rect 191062 227898 191146 228134
rect 191382 227898 226826 228134
rect 227062 227898 227146 228134
rect 227382 227898 262826 228134
rect 263062 227898 263146 228134
rect 263382 227898 298826 228134
rect 299062 227898 299146 228134
rect 299382 227898 334826 228134
rect 335062 227898 335146 228134
rect 335382 227898 370826 228134
rect 371062 227898 371146 228134
rect 371382 227898 406826 228134
rect 407062 227898 407146 228134
rect 407382 227898 442826 228134
rect 443062 227898 443146 228134
rect 443382 227898 478826 228134
rect 479062 227898 479146 228134
rect 479382 227898 514826 228134
rect 515062 227898 515146 228134
rect 515382 227898 550826 228134
rect 551062 227898 551146 228134
rect 551382 227898 587262 228134
rect 587498 227898 587582 228134
rect 587818 227898 592650 228134
rect -8726 227866 592650 227898
rect -8726 223954 592650 223986
rect -8726 223718 -2934 223954
rect -2698 223718 -2614 223954
rect -2378 223718 6326 223954
rect 6562 223718 6646 223954
rect 6882 223718 42326 223954
rect 42562 223718 42646 223954
rect 42882 223718 78326 223954
rect 78562 223718 78646 223954
rect 78882 223718 114326 223954
rect 114562 223718 114646 223954
rect 114882 223718 150326 223954
rect 150562 223718 150646 223954
rect 150882 223718 186326 223954
rect 186562 223718 186646 223954
rect 186882 223718 222326 223954
rect 222562 223718 222646 223954
rect 222882 223718 258326 223954
rect 258562 223718 258646 223954
rect 258882 223718 294326 223954
rect 294562 223718 294646 223954
rect 294882 223718 330326 223954
rect 330562 223718 330646 223954
rect 330882 223718 366326 223954
rect 366562 223718 366646 223954
rect 366882 223718 402326 223954
rect 402562 223718 402646 223954
rect 402882 223718 438326 223954
rect 438562 223718 438646 223954
rect 438882 223718 474326 223954
rect 474562 223718 474646 223954
rect 474882 223718 510326 223954
rect 510562 223718 510646 223954
rect 510882 223718 546326 223954
rect 546562 223718 546646 223954
rect 546882 223718 582326 223954
rect 582562 223718 582646 223954
rect 582882 223718 586302 223954
rect 586538 223718 586622 223954
rect 586858 223718 592650 223954
rect -8726 223634 592650 223718
rect -8726 223398 -2934 223634
rect -2698 223398 -2614 223634
rect -2378 223398 6326 223634
rect 6562 223398 6646 223634
rect 6882 223398 42326 223634
rect 42562 223398 42646 223634
rect 42882 223398 78326 223634
rect 78562 223398 78646 223634
rect 78882 223398 114326 223634
rect 114562 223398 114646 223634
rect 114882 223398 150326 223634
rect 150562 223398 150646 223634
rect 150882 223398 186326 223634
rect 186562 223398 186646 223634
rect 186882 223398 222326 223634
rect 222562 223398 222646 223634
rect 222882 223398 258326 223634
rect 258562 223398 258646 223634
rect 258882 223398 294326 223634
rect 294562 223398 294646 223634
rect 294882 223398 330326 223634
rect 330562 223398 330646 223634
rect 330882 223398 366326 223634
rect 366562 223398 366646 223634
rect 366882 223398 402326 223634
rect 402562 223398 402646 223634
rect 402882 223398 438326 223634
rect 438562 223398 438646 223634
rect 438882 223398 474326 223634
rect 474562 223398 474646 223634
rect 474882 223398 510326 223634
rect 510562 223398 510646 223634
rect 510882 223398 546326 223634
rect 546562 223398 546646 223634
rect 546882 223398 582326 223634
rect 582562 223398 582646 223634
rect 582882 223398 586302 223634
rect 586538 223398 586622 223634
rect 586858 223398 592650 223634
rect -8726 223366 592650 223398
rect -8726 219454 592650 219486
rect -8726 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 592650 219454
rect -8726 219134 592650 219218
rect -8726 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 592650 219134
rect -8726 218866 592650 218898
rect -8726 214954 592650 214986
rect -8726 214718 -8694 214954
rect -8458 214718 -8374 214954
rect -8138 214718 33326 214954
rect 33562 214718 33646 214954
rect 33882 214718 69326 214954
rect 69562 214718 69646 214954
rect 69882 214718 105326 214954
rect 105562 214718 105646 214954
rect 105882 214718 141326 214954
rect 141562 214718 141646 214954
rect 141882 214718 177326 214954
rect 177562 214718 177646 214954
rect 177882 214718 213326 214954
rect 213562 214718 213646 214954
rect 213882 214718 249326 214954
rect 249562 214718 249646 214954
rect 249882 214718 285326 214954
rect 285562 214718 285646 214954
rect 285882 214718 321326 214954
rect 321562 214718 321646 214954
rect 321882 214718 357326 214954
rect 357562 214718 357646 214954
rect 357882 214718 393326 214954
rect 393562 214718 393646 214954
rect 393882 214718 429326 214954
rect 429562 214718 429646 214954
rect 429882 214718 465326 214954
rect 465562 214718 465646 214954
rect 465882 214718 501326 214954
rect 501562 214718 501646 214954
rect 501882 214718 537326 214954
rect 537562 214718 537646 214954
rect 537882 214718 573326 214954
rect 573562 214718 573646 214954
rect 573882 214718 592062 214954
rect 592298 214718 592382 214954
rect 592618 214718 592650 214954
rect -8726 214634 592650 214718
rect -8726 214398 -8694 214634
rect -8458 214398 -8374 214634
rect -8138 214398 33326 214634
rect 33562 214398 33646 214634
rect 33882 214398 69326 214634
rect 69562 214398 69646 214634
rect 69882 214398 105326 214634
rect 105562 214398 105646 214634
rect 105882 214398 141326 214634
rect 141562 214398 141646 214634
rect 141882 214398 177326 214634
rect 177562 214398 177646 214634
rect 177882 214398 213326 214634
rect 213562 214398 213646 214634
rect 213882 214398 249326 214634
rect 249562 214398 249646 214634
rect 249882 214398 285326 214634
rect 285562 214398 285646 214634
rect 285882 214398 321326 214634
rect 321562 214398 321646 214634
rect 321882 214398 357326 214634
rect 357562 214398 357646 214634
rect 357882 214398 393326 214634
rect 393562 214398 393646 214634
rect 393882 214398 429326 214634
rect 429562 214398 429646 214634
rect 429882 214398 465326 214634
rect 465562 214398 465646 214634
rect 465882 214398 501326 214634
rect 501562 214398 501646 214634
rect 501882 214398 537326 214634
rect 537562 214398 537646 214634
rect 537882 214398 573326 214634
rect 573562 214398 573646 214634
rect 573882 214398 592062 214634
rect 592298 214398 592382 214634
rect 592618 214398 592650 214634
rect -8726 214366 592650 214398
rect -8726 210454 592650 210486
rect -8726 210218 -7734 210454
rect -7498 210218 -7414 210454
rect -7178 210218 28826 210454
rect 29062 210218 29146 210454
rect 29382 210218 64826 210454
rect 65062 210218 65146 210454
rect 65382 210218 100826 210454
rect 101062 210218 101146 210454
rect 101382 210218 136826 210454
rect 137062 210218 137146 210454
rect 137382 210218 172826 210454
rect 173062 210218 173146 210454
rect 173382 210218 208826 210454
rect 209062 210218 209146 210454
rect 209382 210218 244826 210454
rect 245062 210218 245146 210454
rect 245382 210218 280826 210454
rect 281062 210218 281146 210454
rect 281382 210218 316826 210454
rect 317062 210218 317146 210454
rect 317382 210218 352826 210454
rect 353062 210218 353146 210454
rect 353382 210218 388826 210454
rect 389062 210218 389146 210454
rect 389382 210218 424826 210454
rect 425062 210218 425146 210454
rect 425382 210218 460826 210454
rect 461062 210218 461146 210454
rect 461382 210218 496826 210454
rect 497062 210218 497146 210454
rect 497382 210218 532826 210454
rect 533062 210218 533146 210454
rect 533382 210218 568826 210454
rect 569062 210218 569146 210454
rect 569382 210218 591102 210454
rect 591338 210218 591422 210454
rect 591658 210218 592650 210454
rect -8726 210134 592650 210218
rect -8726 209898 -7734 210134
rect -7498 209898 -7414 210134
rect -7178 209898 28826 210134
rect 29062 209898 29146 210134
rect 29382 209898 64826 210134
rect 65062 209898 65146 210134
rect 65382 209898 100826 210134
rect 101062 209898 101146 210134
rect 101382 209898 136826 210134
rect 137062 209898 137146 210134
rect 137382 209898 172826 210134
rect 173062 209898 173146 210134
rect 173382 209898 208826 210134
rect 209062 209898 209146 210134
rect 209382 209898 244826 210134
rect 245062 209898 245146 210134
rect 245382 209898 280826 210134
rect 281062 209898 281146 210134
rect 281382 209898 316826 210134
rect 317062 209898 317146 210134
rect 317382 209898 352826 210134
rect 353062 209898 353146 210134
rect 353382 209898 388826 210134
rect 389062 209898 389146 210134
rect 389382 209898 424826 210134
rect 425062 209898 425146 210134
rect 425382 209898 460826 210134
rect 461062 209898 461146 210134
rect 461382 209898 496826 210134
rect 497062 209898 497146 210134
rect 497382 209898 532826 210134
rect 533062 209898 533146 210134
rect 533382 209898 568826 210134
rect 569062 209898 569146 210134
rect 569382 209898 591102 210134
rect 591338 209898 591422 210134
rect 591658 209898 592650 210134
rect -8726 209866 592650 209898
rect -8726 205954 592650 205986
rect -8726 205718 -6774 205954
rect -6538 205718 -6454 205954
rect -6218 205718 24326 205954
rect 24562 205718 24646 205954
rect 24882 205718 60326 205954
rect 60562 205718 60646 205954
rect 60882 205718 96326 205954
rect 96562 205718 96646 205954
rect 96882 205718 132326 205954
rect 132562 205718 132646 205954
rect 132882 205718 168326 205954
rect 168562 205718 168646 205954
rect 168882 205718 204326 205954
rect 204562 205718 204646 205954
rect 204882 205718 240326 205954
rect 240562 205718 240646 205954
rect 240882 205718 276326 205954
rect 276562 205718 276646 205954
rect 276882 205718 312326 205954
rect 312562 205718 312646 205954
rect 312882 205718 348326 205954
rect 348562 205718 348646 205954
rect 348882 205718 384326 205954
rect 384562 205718 384646 205954
rect 384882 205718 420326 205954
rect 420562 205718 420646 205954
rect 420882 205718 456326 205954
rect 456562 205718 456646 205954
rect 456882 205718 492326 205954
rect 492562 205718 492646 205954
rect 492882 205718 528326 205954
rect 528562 205718 528646 205954
rect 528882 205718 564326 205954
rect 564562 205718 564646 205954
rect 564882 205718 590142 205954
rect 590378 205718 590462 205954
rect 590698 205718 592650 205954
rect -8726 205634 592650 205718
rect -8726 205398 -6774 205634
rect -6538 205398 -6454 205634
rect -6218 205398 24326 205634
rect 24562 205398 24646 205634
rect 24882 205398 60326 205634
rect 60562 205398 60646 205634
rect 60882 205398 96326 205634
rect 96562 205398 96646 205634
rect 96882 205398 132326 205634
rect 132562 205398 132646 205634
rect 132882 205398 168326 205634
rect 168562 205398 168646 205634
rect 168882 205398 204326 205634
rect 204562 205398 204646 205634
rect 204882 205398 240326 205634
rect 240562 205398 240646 205634
rect 240882 205398 276326 205634
rect 276562 205398 276646 205634
rect 276882 205398 312326 205634
rect 312562 205398 312646 205634
rect 312882 205398 348326 205634
rect 348562 205398 348646 205634
rect 348882 205398 384326 205634
rect 384562 205398 384646 205634
rect 384882 205398 420326 205634
rect 420562 205398 420646 205634
rect 420882 205398 456326 205634
rect 456562 205398 456646 205634
rect 456882 205398 492326 205634
rect 492562 205398 492646 205634
rect 492882 205398 528326 205634
rect 528562 205398 528646 205634
rect 528882 205398 564326 205634
rect 564562 205398 564646 205634
rect 564882 205398 590142 205634
rect 590378 205398 590462 205634
rect 590698 205398 592650 205634
rect -8726 205366 592650 205398
rect -8726 201454 592650 201486
rect -8726 201218 -5814 201454
rect -5578 201218 -5494 201454
rect -5258 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 127826 201454
rect 128062 201218 128146 201454
rect 128382 201218 163826 201454
rect 164062 201218 164146 201454
rect 164382 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 235826 201454
rect 236062 201218 236146 201454
rect 236382 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 589182 201454
rect 589418 201218 589502 201454
rect 589738 201218 592650 201454
rect -8726 201134 592650 201218
rect -8726 200898 -5814 201134
rect -5578 200898 -5494 201134
rect -5258 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 127826 201134
rect 128062 200898 128146 201134
rect 128382 200898 163826 201134
rect 164062 200898 164146 201134
rect 164382 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 235826 201134
rect 236062 200898 236146 201134
rect 236382 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 589182 201134
rect 589418 200898 589502 201134
rect 589738 200898 592650 201134
rect -8726 200866 592650 200898
rect -8726 196954 592650 196986
rect -8726 196718 -4854 196954
rect -4618 196718 -4534 196954
rect -4298 196718 15326 196954
rect 15562 196718 15646 196954
rect 15882 196718 51326 196954
rect 51562 196718 51646 196954
rect 51882 196718 87326 196954
rect 87562 196718 87646 196954
rect 87882 196718 123326 196954
rect 123562 196718 123646 196954
rect 123882 196718 159326 196954
rect 159562 196718 159646 196954
rect 159882 196718 195326 196954
rect 195562 196718 195646 196954
rect 195882 196718 231326 196954
rect 231562 196718 231646 196954
rect 231882 196718 267326 196954
rect 267562 196718 267646 196954
rect 267882 196718 303326 196954
rect 303562 196718 303646 196954
rect 303882 196718 339326 196954
rect 339562 196718 339646 196954
rect 339882 196718 375326 196954
rect 375562 196718 375646 196954
rect 375882 196718 411326 196954
rect 411562 196718 411646 196954
rect 411882 196718 447326 196954
rect 447562 196718 447646 196954
rect 447882 196718 483326 196954
rect 483562 196718 483646 196954
rect 483882 196718 519326 196954
rect 519562 196718 519646 196954
rect 519882 196718 555326 196954
rect 555562 196718 555646 196954
rect 555882 196718 588222 196954
rect 588458 196718 588542 196954
rect 588778 196718 592650 196954
rect -8726 196634 592650 196718
rect -8726 196398 -4854 196634
rect -4618 196398 -4534 196634
rect -4298 196398 15326 196634
rect 15562 196398 15646 196634
rect 15882 196398 51326 196634
rect 51562 196398 51646 196634
rect 51882 196398 87326 196634
rect 87562 196398 87646 196634
rect 87882 196398 123326 196634
rect 123562 196398 123646 196634
rect 123882 196398 159326 196634
rect 159562 196398 159646 196634
rect 159882 196398 195326 196634
rect 195562 196398 195646 196634
rect 195882 196398 231326 196634
rect 231562 196398 231646 196634
rect 231882 196398 267326 196634
rect 267562 196398 267646 196634
rect 267882 196398 303326 196634
rect 303562 196398 303646 196634
rect 303882 196398 339326 196634
rect 339562 196398 339646 196634
rect 339882 196398 375326 196634
rect 375562 196398 375646 196634
rect 375882 196398 411326 196634
rect 411562 196398 411646 196634
rect 411882 196398 447326 196634
rect 447562 196398 447646 196634
rect 447882 196398 483326 196634
rect 483562 196398 483646 196634
rect 483882 196398 519326 196634
rect 519562 196398 519646 196634
rect 519882 196398 555326 196634
rect 555562 196398 555646 196634
rect 555882 196398 588222 196634
rect 588458 196398 588542 196634
rect 588778 196398 592650 196634
rect -8726 196366 592650 196398
rect -8726 192454 592650 192486
rect -8726 192218 -3894 192454
rect -3658 192218 -3574 192454
rect -3338 192218 10826 192454
rect 11062 192218 11146 192454
rect 11382 192218 46826 192454
rect 47062 192218 47146 192454
rect 47382 192218 82826 192454
rect 83062 192218 83146 192454
rect 83382 192218 118826 192454
rect 119062 192218 119146 192454
rect 119382 192218 154826 192454
rect 155062 192218 155146 192454
rect 155382 192218 190826 192454
rect 191062 192218 191146 192454
rect 191382 192218 226826 192454
rect 227062 192218 227146 192454
rect 227382 192218 262826 192454
rect 263062 192218 263146 192454
rect 263382 192218 298826 192454
rect 299062 192218 299146 192454
rect 299382 192218 334826 192454
rect 335062 192218 335146 192454
rect 335382 192218 370826 192454
rect 371062 192218 371146 192454
rect 371382 192218 406826 192454
rect 407062 192218 407146 192454
rect 407382 192218 442826 192454
rect 443062 192218 443146 192454
rect 443382 192218 478826 192454
rect 479062 192218 479146 192454
rect 479382 192218 514826 192454
rect 515062 192218 515146 192454
rect 515382 192218 550826 192454
rect 551062 192218 551146 192454
rect 551382 192218 587262 192454
rect 587498 192218 587582 192454
rect 587818 192218 592650 192454
rect -8726 192134 592650 192218
rect -8726 191898 -3894 192134
rect -3658 191898 -3574 192134
rect -3338 191898 10826 192134
rect 11062 191898 11146 192134
rect 11382 191898 46826 192134
rect 47062 191898 47146 192134
rect 47382 191898 82826 192134
rect 83062 191898 83146 192134
rect 83382 191898 118826 192134
rect 119062 191898 119146 192134
rect 119382 191898 154826 192134
rect 155062 191898 155146 192134
rect 155382 191898 190826 192134
rect 191062 191898 191146 192134
rect 191382 191898 226826 192134
rect 227062 191898 227146 192134
rect 227382 191898 262826 192134
rect 263062 191898 263146 192134
rect 263382 191898 298826 192134
rect 299062 191898 299146 192134
rect 299382 191898 334826 192134
rect 335062 191898 335146 192134
rect 335382 191898 370826 192134
rect 371062 191898 371146 192134
rect 371382 191898 406826 192134
rect 407062 191898 407146 192134
rect 407382 191898 442826 192134
rect 443062 191898 443146 192134
rect 443382 191898 478826 192134
rect 479062 191898 479146 192134
rect 479382 191898 514826 192134
rect 515062 191898 515146 192134
rect 515382 191898 550826 192134
rect 551062 191898 551146 192134
rect 551382 191898 587262 192134
rect 587498 191898 587582 192134
rect 587818 191898 592650 192134
rect -8726 191866 592650 191898
rect -8726 187954 592650 187986
rect -8726 187718 -2934 187954
rect -2698 187718 -2614 187954
rect -2378 187718 6326 187954
rect 6562 187718 6646 187954
rect 6882 187718 42326 187954
rect 42562 187718 42646 187954
rect 42882 187718 78326 187954
rect 78562 187718 78646 187954
rect 78882 187718 114326 187954
rect 114562 187718 114646 187954
rect 114882 187718 150326 187954
rect 150562 187718 150646 187954
rect 150882 187718 186326 187954
rect 186562 187718 186646 187954
rect 186882 187718 222326 187954
rect 222562 187718 222646 187954
rect 222882 187718 258326 187954
rect 258562 187718 258646 187954
rect 258882 187718 294326 187954
rect 294562 187718 294646 187954
rect 294882 187718 330326 187954
rect 330562 187718 330646 187954
rect 330882 187718 366326 187954
rect 366562 187718 366646 187954
rect 366882 187718 402326 187954
rect 402562 187718 402646 187954
rect 402882 187718 438326 187954
rect 438562 187718 438646 187954
rect 438882 187718 474326 187954
rect 474562 187718 474646 187954
rect 474882 187718 510326 187954
rect 510562 187718 510646 187954
rect 510882 187718 546326 187954
rect 546562 187718 546646 187954
rect 546882 187718 582326 187954
rect 582562 187718 582646 187954
rect 582882 187718 586302 187954
rect 586538 187718 586622 187954
rect 586858 187718 592650 187954
rect -8726 187634 592650 187718
rect -8726 187398 -2934 187634
rect -2698 187398 -2614 187634
rect -2378 187398 6326 187634
rect 6562 187398 6646 187634
rect 6882 187398 42326 187634
rect 42562 187398 42646 187634
rect 42882 187398 78326 187634
rect 78562 187398 78646 187634
rect 78882 187398 114326 187634
rect 114562 187398 114646 187634
rect 114882 187398 150326 187634
rect 150562 187398 150646 187634
rect 150882 187398 186326 187634
rect 186562 187398 186646 187634
rect 186882 187398 222326 187634
rect 222562 187398 222646 187634
rect 222882 187398 258326 187634
rect 258562 187398 258646 187634
rect 258882 187398 294326 187634
rect 294562 187398 294646 187634
rect 294882 187398 330326 187634
rect 330562 187398 330646 187634
rect 330882 187398 366326 187634
rect 366562 187398 366646 187634
rect 366882 187398 402326 187634
rect 402562 187398 402646 187634
rect 402882 187398 438326 187634
rect 438562 187398 438646 187634
rect 438882 187398 474326 187634
rect 474562 187398 474646 187634
rect 474882 187398 510326 187634
rect 510562 187398 510646 187634
rect 510882 187398 546326 187634
rect 546562 187398 546646 187634
rect 546882 187398 582326 187634
rect 582562 187398 582646 187634
rect 582882 187398 586302 187634
rect 586538 187398 586622 187634
rect 586858 187398 592650 187634
rect -8726 187366 592650 187398
rect -8726 183454 592650 183486
rect -8726 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 592650 183454
rect -8726 183134 592650 183218
rect -8726 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 592650 183134
rect -8726 182866 592650 182898
rect -8726 178954 592650 178986
rect -8726 178718 -8694 178954
rect -8458 178718 -8374 178954
rect -8138 178718 33326 178954
rect 33562 178718 33646 178954
rect 33882 178718 69326 178954
rect 69562 178718 69646 178954
rect 69882 178718 105326 178954
rect 105562 178718 105646 178954
rect 105882 178718 141326 178954
rect 141562 178718 141646 178954
rect 141882 178718 177326 178954
rect 177562 178718 177646 178954
rect 177882 178718 213326 178954
rect 213562 178718 213646 178954
rect 213882 178718 249326 178954
rect 249562 178718 249646 178954
rect 249882 178718 285326 178954
rect 285562 178718 285646 178954
rect 285882 178718 321326 178954
rect 321562 178718 321646 178954
rect 321882 178718 357326 178954
rect 357562 178718 357646 178954
rect 357882 178718 393326 178954
rect 393562 178718 393646 178954
rect 393882 178718 429326 178954
rect 429562 178718 429646 178954
rect 429882 178718 465326 178954
rect 465562 178718 465646 178954
rect 465882 178718 501326 178954
rect 501562 178718 501646 178954
rect 501882 178718 537326 178954
rect 537562 178718 537646 178954
rect 537882 178718 573326 178954
rect 573562 178718 573646 178954
rect 573882 178718 592062 178954
rect 592298 178718 592382 178954
rect 592618 178718 592650 178954
rect -8726 178634 592650 178718
rect -8726 178398 -8694 178634
rect -8458 178398 -8374 178634
rect -8138 178398 33326 178634
rect 33562 178398 33646 178634
rect 33882 178398 69326 178634
rect 69562 178398 69646 178634
rect 69882 178398 105326 178634
rect 105562 178398 105646 178634
rect 105882 178398 141326 178634
rect 141562 178398 141646 178634
rect 141882 178398 177326 178634
rect 177562 178398 177646 178634
rect 177882 178398 213326 178634
rect 213562 178398 213646 178634
rect 213882 178398 249326 178634
rect 249562 178398 249646 178634
rect 249882 178398 285326 178634
rect 285562 178398 285646 178634
rect 285882 178398 321326 178634
rect 321562 178398 321646 178634
rect 321882 178398 357326 178634
rect 357562 178398 357646 178634
rect 357882 178398 393326 178634
rect 393562 178398 393646 178634
rect 393882 178398 429326 178634
rect 429562 178398 429646 178634
rect 429882 178398 465326 178634
rect 465562 178398 465646 178634
rect 465882 178398 501326 178634
rect 501562 178398 501646 178634
rect 501882 178398 537326 178634
rect 537562 178398 537646 178634
rect 537882 178398 573326 178634
rect 573562 178398 573646 178634
rect 573882 178398 592062 178634
rect 592298 178398 592382 178634
rect 592618 178398 592650 178634
rect -8726 178366 592650 178398
rect -8726 174454 592650 174486
rect -8726 174218 -7734 174454
rect -7498 174218 -7414 174454
rect -7178 174218 28826 174454
rect 29062 174218 29146 174454
rect 29382 174218 64826 174454
rect 65062 174218 65146 174454
rect 65382 174218 100826 174454
rect 101062 174218 101146 174454
rect 101382 174218 136826 174454
rect 137062 174218 137146 174454
rect 137382 174218 172826 174454
rect 173062 174218 173146 174454
rect 173382 174218 208826 174454
rect 209062 174218 209146 174454
rect 209382 174218 244826 174454
rect 245062 174218 245146 174454
rect 245382 174218 280826 174454
rect 281062 174218 281146 174454
rect 281382 174218 316826 174454
rect 317062 174218 317146 174454
rect 317382 174218 352826 174454
rect 353062 174218 353146 174454
rect 353382 174218 388826 174454
rect 389062 174218 389146 174454
rect 389382 174218 424826 174454
rect 425062 174218 425146 174454
rect 425382 174218 460826 174454
rect 461062 174218 461146 174454
rect 461382 174218 496826 174454
rect 497062 174218 497146 174454
rect 497382 174218 532826 174454
rect 533062 174218 533146 174454
rect 533382 174218 568826 174454
rect 569062 174218 569146 174454
rect 569382 174218 591102 174454
rect 591338 174218 591422 174454
rect 591658 174218 592650 174454
rect -8726 174134 592650 174218
rect -8726 173898 -7734 174134
rect -7498 173898 -7414 174134
rect -7178 173898 28826 174134
rect 29062 173898 29146 174134
rect 29382 173898 64826 174134
rect 65062 173898 65146 174134
rect 65382 173898 100826 174134
rect 101062 173898 101146 174134
rect 101382 173898 136826 174134
rect 137062 173898 137146 174134
rect 137382 173898 172826 174134
rect 173062 173898 173146 174134
rect 173382 173898 208826 174134
rect 209062 173898 209146 174134
rect 209382 173898 244826 174134
rect 245062 173898 245146 174134
rect 245382 173898 280826 174134
rect 281062 173898 281146 174134
rect 281382 173898 316826 174134
rect 317062 173898 317146 174134
rect 317382 173898 352826 174134
rect 353062 173898 353146 174134
rect 353382 173898 388826 174134
rect 389062 173898 389146 174134
rect 389382 173898 424826 174134
rect 425062 173898 425146 174134
rect 425382 173898 460826 174134
rect 461062 173898 461146 174134
rect 461382 173898 496826 174134
rect 497062 173898 497146 174134
rect 497382 173898 532826 174134
rect 533062 173898 533146 174134
rect 533382 173898 568826 174134
rect 569062 173898 569146 174134
rect 569382 173898 591102 174134
rect 591338 173898 591422 174134
rect 591658 173898 592650 174134
rect -8726 173866 592650 173898
rect -8726 169954 592650 169986
rect -8726 169718 -6774 169954
rect -6538 169718 -6454 169954
rect -6218 169718 24326 169954
rect 24562 169718 24646 169954
rect 24882 169718 60326 169954
rect 60562 169718 60646 169954
rect 60882 169718 96326 169954
rect 96562 169718 96646 169954
rect 96882 169718 132326 169954
rect 132562 169718 132646 169954
rect 132882 169718 168326 169954
rect 168562 169718 168646 169954
rect 168882 169718 204326 169954
rect 204562 169718 204646 169954
rect 204882 169718 240326 169954
rect 240562 169718 240646 169954
rect 240882 169718 276326 169954
rect 276562 169718 276646 169954
rect 276882 169718 312326 169954
rect 312562 169718 312646 169954
rect 312882 169718 348326 169954
rect 348562 169718 348646 169954
rect 348882 169718 384326 169954
rect 384562 169718 384646 169954
rect 384882 169718 420326 169954
rect 420562 169718 420646 169954
rect 420882 169718 456326 169954
rect 456562 169718 456646 169954
rect 456882 169718 492326 169954
rect 492562 169718 492646 169954
rect 492882 169718 528326 169954
rect 528562 169718 528646 169954
rect 528882 169718 564326 169954
rect 564562 169718 564646 169954
rect 564882 169718 590142 169954
rect 590378 169718 590462 169954
rect 590698 169718 592650 169954
rect -8726 169634 592650 169718
rect -8726 169398 -6774 169634
rect -6538 169398 -6454 169634
rect -6218 169398 24326 169634
rect 24562 169398 24646 169634
rect 24882 169398 60326 169634
rect 60562 169398 60646 169634
rect 60882 169398 96326 169634
rect 96562 169398 96646 169634
rect 96882 169398 132326 169634
rect 132562 169398 132646 169634
rect 132882 169398 168326 169634
rect 168562 169398 168646 169634
rect 168882 169398 204326 169634
rect 204562 169398 204646 169634
rect 204882 169398 240326 169634
rect 240562 169398 240646 169634
rect 240882 169398 276326 169634
rect 276562 169398 276646 169634
rect 276882 169398 312326 169634
rect 312562 169398 312646 169634
rect 312882 169398 348326 169634
rect 348562 169398 348646 169634
rect 348882 169398 384326 169634
rect 384562 169398 384646 169634
rect 384882 169398 420326 169634
rect 420562 169398 420646 169634
rect 420882 169398 456326 169634
rect 456562 169398 456646 169634
rect 456882 169398 492326 169634
rect 492562 169398 492646 169634
rect 492882 169398 528326 169634
rect 528562 169398 528646 169634
rect 528882 169398 564326 169634
rect 564562 169398 564646 169634
rect 564882 169398 590142 169634
rect 590378 169398 590462 169634
rect 590698 169398 592650 169634
rect -8726 169366 592650 169398
rect -8726 165454 592650 165486
rect -8726 165218 -5814 165454
rect -5578 165218 -5494 165454
rect -5258 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 91826 165454
rect 92062 165218 92146 165454
rect 92382 165218 127826 165454
rect 128062 165218 128146 165454
rect 128382 165218 163826 165454
rect 164062 165218 164146 165454
rect 164382 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 235826 165454
rect 236062 165218 236146 165454
rect 236382 165218 271826 165454
rect 272062 165218 272146 165454
rect 272382 165218 307826 165454
rect 308062 165218 308146 165454
rect 308382 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 589182 165454
rect 589418 165218 589502 165454
rect 589738 165218 592650 165454
rect -8726 165134 592650 165218
rect -8726 164898 -5814 165134
rect -5578 164898 -5494 165134
rect -5258 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 91826 165134
rect 92062 164898 92146 165134
rect 92382 164898 127826 165134
rect 128062 164898 128146 165134
rect 128382 164898 163826 165134
rect 164062 164898 164146 165134
rect 164382 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 235826 165134
rect 236062 164898 236146 165134
rect 236382 164898 271826 165134
rect 272062 164898 272146 165134
rect 272382 164898 307826 165134
rect 308062 164898 308146 165134
rect 308382 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 589182 165134
rect 589418 164898 589502 165134
rect 589738 164898 592650 165134
rect -8726 164866 592650 164898
rect -8726 160954 592650 160986
rect -8726 160718 -4854 160954
rect -4618 160718 -4534 160954
rect -4298 160718 15326 160954
rect 15562 160718 15646 160954
rect 15882 160718 51326 160954
rect 51562 160718 51646 160954
rect 51882 160718 87326 160954
rect 87562 160718 87646 160954
rect 87882 160718 123326 160954
rect 123562 160718 123646 160954
rect 123882 160718 159326 160954
rect 159562 160718 159646 160954
rect 159882 160718 195326 160954
rect 195562 160718 195646 160954
rect 195882 160718 231326 160954
rect 231562 160718 231646 160954
rect 231882 160718 267326 160954
rect 267562 160718 267646 160954
rect 267882 160718 303326 160954
rect 303562 160718 303646 160954
rect 303882 160718 339326 160954
rect 339562 160718 339646 160954
rect 339882 160718 375326 160954
rect 375562 160718 375646 160954
rect 375882 160718 411326 160954
rect 411562 160718 411646 160954
rect 411882 160718 447326 160954
rect 447562 160718 447646 160954
rect 447882 160718 483326 160954
rect 483562 160718 483646 160954
rect 483882 160718 519326 160954
rect 519562 160718 519646 160954
rect 519882 160718 555326 160954
rect 555562 160718 555646 160954
rect 555882 160718 588222 160954
rect 588458 160718 588542 160954
rect 588778 160718 592650 160954
rect -8726 160634 592650 160718
rect -8726 160398 -4854 160634
rect -4618 160398 -4534 160634
rect -4298 160398 15326 160634
rect 15562 160398 15646 160634
rect 15882 160398 51326 160634
rect 51562 160398 51646 160634
rect 51882 160398 87326 160634
rect 87562 160398 87646 160634
rect 87882 160398 123326 160634
rect 123562 160398 123646 160634
rect 123882 160398 159326 160634
rect 159562 160398 159646 160634
rect 159882 160398 195326 160634
rect 195562 160398 195646 160634
rect 195882 160398 231326 160634
rect 231562 160398 231646 160634
rect 231882 160398 267326 160634
rect 267562 160398 267646 160634
rect 267882 160398 303326 160634
rect 303562 160398 303646 160634
rect 303882 160398 339326 160634
rect 339562 160398 339646 160634
rect 339882 160398 375326 160634
rect 375562 160398 375646 160634
rect 375882 160398 411326 160634
rect 411562 160398 411646 160634
rect 411882 160398 447326 160634
rect 447562 160398 447646 160634
rect 447882 160398 483326 160634
rect 483562 160398 483646 160634
rect 483882 160398 519326 160634
rect 519562 160398 519646 160634
rect 519882 160398 555326 160634
rect 555562 160398 555646 160634
rect 555882 160398 588222 160634
rect 588458 160398 588542 160634
rect 588778 160398 592650 160634
rect -8726 160366 592650 160398
rect -8726 156454 592650 156486
rect -8726 156218 -3894 156454
rect -3658 156218 -3574 156454
rect -3338 156218 10826 156454
rect 11062 156218 11146 156454
rect 11382 156218 46826 156454
rect 47062 156218 47146 156454
rect 47382 156218 82826 156454
rect 83062 156218 83146 156454
rect 83382 156218 118826 156454
rect 119062 156218 119146 156454
rect 119382 156218 154826 156454
rect 155062 156218 155146 156454
rect 155382 156218 190826 156454
rect 191062 156218 191146 156454
rect 191382 156218 226826 156454
rect 227062 156218 227146 156454
rect 227382 156218 370826 156454
rect 371062 156218 371146 156454
rect 371382 156218 406826 156454
rect 407062 156218 407146 156454
rect 407382 156218 442826 156454
rect 443062 156218 443146 156454
rect 443382 156218 478826 156454
rect 479062 156218 479146 156454
rect 479382 156218 514826 156454
rect 515062 156218 515146 156454
rect 515382 156218 550826 156454
rect 551062 156218 551146 156454
rect 551382 156218 587262 156454
rect 587498 156218 587582 156454
rect 587818 156218 592650 156454
rect -8726 156134 592650 156218
rect -8726 155898 -3894 156134
rect -3658 155898 -3574 156134
rect -3338 155898 10826 156134
rect 11062 155898 11146 156134
rect 11382 155898 46826 156134
rect 47062 155898 47146 156134
rect 47382 155898 82826 156134
rect 83062 155898 83146 156134
rect 83382 155898 118826 156134
rect 119062 155898 119146 156134
rect 119382 155898 154826 156134
rect 155062 155898 155146 156134
rect 155382 155898 190826 156134
rect 191062 155898 191146 156134
rect 191382 155898 226826 156134
rect 227062 155898 227146 156134
rect 227382 155898 370826 156134
rect 371062 155898 371146 156134
rect 371382 155898 406826 156134
rect 407062 155898 407146 156134
rect 407382 155898 442826 156134
rect 443062 155898 443146 156134
rect 443382 155898 478826 156134
rect 479062 155898 479146 156134
rect 479382 155898 514826 156134
rect 515062 155898 515146 156134
rect 515382 155898 550826 156134
rect 551062 155898 551146 156134
rect 551382 155898 587262 156134
rect 587498 155898 587582 156134
rect 587818 155898 592650 156134
rect -8726 155866 592650 155898
rect -8726 151954 592650 151986
rect -8726 151718 -2934 151954
rect -2698 151718 -2614 151954
rect -2378 151718 6326 151954
rect 6562 151718 6646 151954
rect 6882 151718 42326 151954
rect 42562 151718 42646 151954
rect 42882 151718 78326 151954
rect 78562 151718 78646 151954
rect 78882 151718 114326 151954
rect 114562 151718 114646 151954
rect 114882 151718 150326 151954
rect 150562 151718 150646 151954
rect 150882 151718 186326 151954
rect 186562 151718 186646 151954
rect 186882 151718 222326 151954
rect 222562 151718 222646 151954
rect 222882 151718 279610 151954
rect 279846 151718 310330 151954
rect 310566 151718 341050 151954
rect 341286 151718 366326 151954
rect 366562 151718 366646 151954
rect 366882 151718 402326 151954
rect 402562 151718 402646 151954
rect 402882 151718 438326 151954
rect 438562 151718 438646 151954
rect 438882 151718 474326 151954
rect 474562 151718 474646 151954
rect 474882 151718 510326 151954
rect 510562 151718 510646 151954
rect 510882 151718 546326 151954
rect 546562 151718 546646 151954
rect 546882 151718 582326 151954
rect 582562 151718 582646 151954
rect 582882 151718 586302 151954
rect 586538 151718 586622 151954
rect 586858 151718 592650 151954
rect -8726 151634 592650 151718
rect -8726 151398 -2934 151634
rect -2698 151398 -2614 151634
rect -2378 151398 6326 151634
rect 6562 151398 6646 151634
rect 6882 151398 42326 151634
rect 42562 151398 42646 151634
rect 42882 151398 78326 151634
rect 78562 151398 78646 151634
rect 78882 151398 114326 151634
rect 114562 151398 114646 151634
rect 114882 151398 150326 151634
rect 150562 151398 150646 151634
rect 150882 151398 186326 151634
rect 186562 151398 186646 151634
rect 186882 151398 222326 151634
rect 222562 151398 222646 151634
rect 222882 151398 279610 151634
rect 279846 151398 310330 151634
rect 310566 151398 341050 151634
rect 341286 151398 366326 151634
rect 366562 151398 366646 151634
rect 366882 151398 402326 151634
rect 402562 151398 402646 151634
rect 402882 151398 438326 151634
rect 438562 151398 438646 151634
rect 438882 151398 474326 151634
rect 474562 151398 474646 151634
rect 474882 151398 510326 151634
rect 510562 151398 510646 151634
rect 510882 151398 546326 151634
rect 546562 151398 546646 151634
rect 546882 151398 582326 151634
rect 582562 151398 582646 151634
rect 582882 151398 586302 151634
rect 586538 151398 586622 151634
rect 586858 151398 592650 151634
rect -8726 151366 592650 151398
rect -8726 147454 592650 147486
rect -8726 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 264250 147454
rect 264486 147218 294970 147454
rect 295206 147218 325690 147454
rect 325926 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 592650 147454
rect -8726 147134 592650 147218
rect -8726 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 264250 147134
rect 264486 146898 294970 147134
rect 295206 146898 325690 147134
rect 325926 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 592650 147134
rect -8726 146866 592650 146898
rect -8726 142954 592650 142986
rect -8726 142718 -8694 142954
rect -8458 142718 -8374 142954
rect -8138 142718 33326 142954
rect 33562 142718 33646 142954
rect 33882 142718 69326 142954
rect 69562 142718 69646 142954
rect 69882 142718 105326 142954
rect 105562 142718 105646 142954
rect 105882 142718 141326 142954
rect 141562 142718 141646 142954
rect 141882 142718 177326 142954
rect 177562 142718 177646 142954
rect 177882 142718 213326 142954
rect 213562 142718 213646 142954
rect 213882 142718 249326 142954
rect 249562 142718 249646 142954
rect 249882 142718 357326 142954
rect 357562 142718 357646 142954
rect 357882 142718 393326 142954
rect 393562 142718 393646 142954
rect 393882 142718 429326 142954
rect 429562 142718 429646 142954
rect 429882 142718 465326 142954
rect 465562 142718 465646 142954
rect 465882 142718 501326 142954
rect 501562 142718 501646 142954
rect 501882 142718 537326 142954
rect 537562 142718 537646 142954
rect 537882 142718 573326 142954
rect 573562 142718 573646 142954
rect 573882 142718 592062 142954
rect 592298 142718 592382 142954
rect 592618 142718 592650 142954
rect -8726 142634 592650 142718
rect -8726 142398 -8694 142634
rect -8458 142398 -8374 142634
rect -8138 142398 33326 142634
rect 33562 142398 33646 142634
rect 33882 142398 69326 142634
rect 69562 142398 69646 142634
rect 69882 142398 105326 142634
rect 105562 142398 105646 142634
rect 105882 142398 141326 142634
rect 141562 142398 141646 142634
rect 141882 142398 177326 142634
rect 177562 142398 177646 142634
rect 177882 142398 213326 142634
rect 213562 142398 213646 142634
rect 213882 142398 249326 142634
rect 249562 142398 249646 142634
rect 249882 142398 357326 142634
rect 357562 142398 357646 142634
rect 357882 142398 393326 142634
rect 393562 142398 393646 142634
rect 393882 142398 429326 142634
rect 429562 142398 429646 142634
rect 429882 142398 465326 142634
rect 465562 142398 465646 142634
rect 465882 142398 501326 142634
rect 501562 142398 501646 142634
rect 501882 142398 537326 142634
rect 537562 142398 537646 142634
rect 537882 142398 573326 142634
rect 573562 142398 573646 142634
rect 573882 142398 592062 142634
rect 592298 142398 592382 142634
rect 592618 142398 592650 142634
rect -8726 142366 592650 142398
rect -8726 138454 592650 138486
rect -8726 138218 -7734 138454
rect -7498 138218 -7414 138454
rect -7178 138218 28826 138454
rect 29062 138218 29146 138454
rect 29382 138218 64826 138454
rect 65062 138218 65146 138454
rect 65382 138218 100826 138454
rect 101062 138218 101146 138454
rect 101382 138218 136826 138454
rect 137062 138218 137146 138454
rect 137382 138218 172826 138454
rect 173062 138218 173146 138454
rect 173382 138218 208826 138454
rect 209062 138218 209146 138454
rect 209382 138218 244826 138454
rect 245062 138218 245146 138454
rect 245382 138218 352826 138454
rect 353062 138218 353146 138454
rect 353382 138218 388826 138454
rect 389062 138218 389146 138454
rect 389382 138218 424826 138454
rect 425062 138218 425146 138454
rect 425382 138218 460826 138454
rect 461062 138218 461146 138454
rect 461382 138218 496826 138454
rect 497062 138218 497146 138454
rect 497382 138218 532826 138454
rect 533062 138218 533146 138454
rect 533382 138218 568826 138454
rect 569062 138218 569146 138454
rect 569382 138218 591102 138454
rect 591338 138218 591422 138454
rect 591658 138218 592650 138454
rect -8726 138134 592650 138218
rect -8726 137898 -7734 138134
rect -7498 137898 -7414 138134
rect -7178 137898 28826 138134
rect 29062 137898 29146 138134
rect 29382 137898 64826 138134
rect 65062 137898 65146 138134
rect 65382 137898 100826 138134
rect 101062 137898 101146 138134
rect 101382 137898 136826 138134
rect 137062 137898 137146 138134
rect 137382 137898 172826 138134
rect 173062 137898 173146 138134
rect 173382 137898 208826 138134
rect 209062 137898 209146 138134
rect 209382 137898 244826 138134
rect 245062 137898 245146 138134
rect 245382 137898 352826 138134
rect 353062 137898 353146 138134
rect 353382 137898 388826 138134
rect 389062 137898 389146 138134
rect 389382 137898 424826 138134
rect 425062 137898 425146 138134
rect 425382 137898 460826 138134
rect 461062 137898 461146 138134
rect 461382 137898 496826 138134
rect 497062 137898 497146 138134
rect 497382 137898 532826 138134
rect 533062 137898 533146 138134
rect 533382 137898 568826 138134
rect 569062 137898 569146 138134
rect 569382 137898 591102 138134
rect 591338 137898 591422 138134
rect 591658 137898 592650 138134
rect -8726 137866 592650 137898
rect -8726 133954 592650 133986
rect -8726 133718 -6774 133954
rect -6538 133718 -6454 133954
rect -6218 133718 24326 133954
rect 24562 133718 24646 133954
rect 24882 133718 60326 133954
rect 60562 133718 60646 133954
rect 60882 133718 96326 133954
rect 96562 133718 96646 133954
rect 96882 133718 132326 133954
rect 132562 133718 132646 133954
rect 132882 133718 168326 133954
rect 168562 133718 168646 133954
rect 168882 133718 204326 133954
rect 204562 133718 204646 133954
rect 204882 133718 240326 133954
rect 240562 133718 240646 133954
rect 240882 133718 348326 133954
rect 348562 133718 348646 133954
rect 348882 133718 384326 133954
rect 384562 133718 384646 133954
rect 384882 133718 420326 133954
rect 420562 133718 420646 133954
rect 420882 133718 456326 133954
rect 456562 133718 456646 133954
rect 456882 133718 492326 133954
rect 492562 133718 492646 133954
rect 492882 133718 528326 133954
rect 528562 133718 528646 133954
rect 528882 133718 564326 133954
rect 564562 133718 564646 133954
rect 564882 133718 590142 133954
rect 590378 133718 590462 133954
rect 590698 133718 592650 133954
rect -8726 133634 592650 133718
rect -8726 133398 -6774 133634
rect -6538 133398 -6454 133634
rect -6218 133398 24326 133634
rect 24562 133398 24646 133634
rect 24882 133398 60326 133634
rect 60562 133398 60646 133634
rect 60882 133398 96326 133634
rect 96562 133398 96646 133634
rect 96882 133398 132326 133634
rect 132562 133398 132646 133634
rect 132882 133398 168326 133634
rect 168562 133398 168646 133634
rect 168882 133398 204326 133634
rect 204562 133398 204646 133634
rect 204882 133398 240326 133634
rect 240562 133398 240646 133634
rect 240882 133398 348326 133634
rect 348562 133398 348646 133634
rect 348882 133398 384326 133634
rect 384562 133398 384646 133634
rect 384882 133398 420326 133634
rect 420562 133398 420646 133634
rect 420882 133398 456326 133634
rect 456562 133398 456646 133634
rect 456882 133398 492326 133634
rect 492562 133398 492646 133634
rect 492882 133398 528326 133634
rect 528562 133398 528646 133634
rect 528882 133398 564326 133634
rect 564562 133398 564646 133634
rect 564882 133398 590142 133634
rect 590378 133398 590462 133634
rect 590698 133398 592650 133634
rect -8726 133366 592650 133398
rect -8726 129454 592650 129486
rect -8726 129218 -5814 129454
rect -5578 129218 -5494 129454
rect -5258 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 91826 129454
rect 92062 129218 92146 129454
rect 92382 129218 127826 129454
rect 128062 129218 128146 129454
rect 128382 129218 163826 129454
rect 164062 129218 164146 129454
rect 164382 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 589182 129454
rect 589418 129218 589502 129454
rect 589738 129218 592650 129454
rect -8726 129134 592650 129218
rect -8726 128898 -5814 129134
rect -5578 128898 -5494 129134
rect -5258 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 91826 129134
rect 92062 128898 92146 129134
rect 92382 128898 127826 129134
rect 128062 128898 128146 129134
rect 128382 128898 163826 129134
rect 164062 128898 164146 129134
rect 164382 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 589182 129134
rect 589418 128898 589502 129134
rect 589738 128898 592650 129134
rect -8726 128866 592650 128898
rect -8726 124954 592650 124986
rect -8726 124718 -4854 124954
rect -4618 124718 -4534 124954
rect -4298 124718 15326 124954
rect 15562 124718 15646 124954
rect 15882 124718 51326 124954
rect 51562 124718 51646 124954
rect 51882 124718 87326 124954
rect 87562 124718 87646 124954
rect 87882 124718 123326 124954
rect 123562 124718 123646 124954
rect 123882 124718 159326 124954
rect 159562 124718 159646 124954
rect 159882 124718 195326 124954
rect 195562 124718 195646 124954
rect 195882 124718 231326 124954
rect 231562 124718 231646 124954
rect 231882 124718 375326 124954
rect 375562 124718 375646 124954
rect 375882 124718 411326 124954
rect 411562 124718 411646 124954
rect 411882 124718 447326 124954
rect 447562 124718 447646 124954
rect 447882 124718 483326 124954
rect 483562 124718 483646 124954
rect 483882 124718 519326 124954
rect 519562 124718 519646 124954
rect 519882 124718 555326 124954
rect 555562 124718 555646 124954
rect 555882 124718 588222 124954
rect 588458 124718 588542 124954
rect 588778 124718 592650 124954
rect -8726 124634 592650 124718
rect -8726 124398 -4854 124634
rect -4618 124398 -4534 124634
rect -4298 124398 15326 124634
rect 15562 124398 15646 124634
rect 15882 124398 51326 124634
rect 51562 124398 51646 124634
rect 51882 124398 87326 124634
rect 87562 124398 87646 124634
rect 87882 124398 123326 124634
rect 123562 124398 123646 124634
rect 123882 124398 159326 124634
rect 159562 124398 159646 124634
rect 159882 124398 195326 124634
rect 195562 124398 195646 124634
rect 195882 124398 231326 124634
rect 231562 124398 231646 124634
rect 231882 124398 375326 124634
rect 375562 124398 375646 124634
rect 375882 124398 411326 124634
rect 411562 124398 411646 124634
rect 411882 124398 447326 124634
rect 447562 124398 447646 124634
rect 447882 124398 483326 124634
rect 483562 124398 483646 124634
rect 483882 124398 519326 124634
rect 519562 124398 519646 124634
rect 519882 124398 555326 124634
rect 555562 124398 555646 124634
rect 555882 124398 588222 124634
rect 588458 124398 588542 124634
rect 588778 124398 592650 124634
rect -8726 124366 592650 124398
rect -8726 120454 592650 120486
rect -8726 120218 -3894 120454
rect -3658 120218 -3574 120454
rect -3338 120218 10826 120454
rect 11062 120218 11146 120454
rect 11382 120218 46826 120454
rect 47062 120218 47146 120454
rect 47382 120218 82826 120454
rect 83062 120218 83146 120454
rect 83382 120218 118826 120454
rect 119062 120218 119146 120454
rect 119382 120218 154826 120454
rect 155062 120218 155146 120454
rect 155382 120218 190826 120454
rect 191062 120218 191146 120454
rect 191382 120218 226826 120454
rect 227062 120218 227146 120454
rect 227382 120218 370826 120454
rect 371062 120218 371146 120454
rect 371382 120218 406826 120454
rect 407062 120218 407146 120454
rect 407382 120218 442826 120454
rect 443062 120218 443146 120454
rect 443382 120218 478826 120454
rect 479062 120218 479146 120454
rect 479382 120218 514826 120454
rect 515062 120218 515146 120454
rect 515382 120218 550826 120454
rect 551062 120218 551146 120454
rect 551382 120218 587262 120454
rect 587498 120218 587582 120454
rect 587818 120218 592650 120454
rect -8726 120134 592650 120218
rect -8726 119898 -3894 120134
rect -3658 119898 -3574 120134
rect -3338 119898 10826 120134
rect 11062 119898 11146 120134
rect 11382 119898 46826 120134
rect 47062 119898 47146 120134
rect 47382 119898 82826 120134
rect 83062 119898 83146 120134
rect 83382 119898 118826 120134
rect 119062 119898 119146 120134
rect 119382 119898 154826 120134
rect 155062 119898 155146 120134
rect 155382 119898 190826 120134
rect 191062 119898 191146 120134
rect 191382 119898 226826 120134
rect 227062 119898 227146 120134
rect 227382 119898 370826 120134
rect 371062 119898 371146 120134
rect 371382 119898 406826 120134
rect 407062 119898 407146 120134
rect 407382 119898 442826 120134
rect 443062 119898 443146 120134
rect 443382 119898 478826 120134
rect 479062 119898 479146 120134
rect 479382 119898 514826 120134
rect 515062 119898 515146 120134
rect 515382 119898 550826 120134
rect 551062 119898 551146 120134
rect 551382 119898 587262 120134
rect 587498 119898 587582 120134
rect 587818 119898 592650 120134
rect -8726 119866 592650 119898
rect -8726 115954 592650 115986
rect -8726 115718 -2934 115954
rect -2698 115718 -2614 115954
rect -2378 115718 6326 115954
rect 6562 115718 6646 115954
rect 6882 115718 42326 115954
rect 42562 115718 42646 115954
rect 42882 115718 78326 115954
rect 78562 115718 78646 115954
rect 78882 115718 114326 115954
rect 114562 115718 114646 115954
rect 114882 115718 150326 115954
rect 150562 115718 150646 115954
rect 150882 115718 186326 115954
rect 186562 115718 186646 115954
rect 186882 115718 222326 115954
rect 222562 115718 222646 115954
rect 222882 115718 279610 115954
rect 279846 115718 310330 115954
rect 310566 115718 341050 115954
rect 341286 115718 366326 115954
rect 366562 115718 366646 115954
rect 366882 115718 402326 115954
rect 402562 115718 402646 115954
rect 402882 115718 438326 115954
rect 438562 115718 438646 115954
rect 438882 115718 474326 115954
rect 474562 115718 474646 115954
rect 474882 115718 510326 115954
rect 510562 115718 510646 115954
rect 510882 115718 546326 115954
rect 546562 115718 546646 115954
rect 546882 115718 582326 115954
rect 582562 115718 582646 115954
rect 582882 115718 586302 115954
rect 586538 115718 586622 115954
rect 586858 115718 592650 115954
rect -8726 115634 592650 115718
rect -8726 115398 -2934 115634
rect -2698 115398 -2614 115634
rect -2378 115398 6326 115634
rect 6562 115398 6646 115634
rect 6882 115398 42326 115634
rect 42562 115398 42646 115634
rect 42882 115398 78326 115634
rect 78562 115398 78646 115634
rect 78882 115398 114326 115634
rect 114562 115398 114646 115634
rect 114882 115398 150326 115634
rect 150562 115398 150646 115634
rect 150882 115398 186326 115634
rect 186562 115398 186646 115634
rect 186882 115398 222326 115634
rect 222562 115398 222646 115634
rect 222882 115398 279610 115634
rect 279846 115398 310330 115634
rect 310566 115398 341050 115634
rect 341286 115398 366326 115634
rect 366562 115398 366646 115634
rect 366882 115398 402326 115634
rect 402562 115398 402646 115634
rect 402882 115398 438326 115634
rect 438562 115398 438646 115634
rect 438882 115398 474326 115634
rect 474562 115398 474646 115634
rect 474882 115398 510326 115634
rect 510562 115398 510646 115634
rect 510882 115398 546326 115634
rect 546562 115398 546646 115634
rect 546882 115398 582326 115634
rect 582562 115398 582646 115634
rect 582882 115398 586302 115634
rect 586538 115398 586622 115634
rect 586858 115398 592650 115634
rect -8726 115366 592650 115398
rect -8726 111454 592650 111486
rect -8726 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 73826 111454
rect 74062 111218 74146 111454
rect 74382 111218 109826 111454
rect 110062 111218 110146 111454
rect 110382 111218 145826 111454
rect 146062 111218 146146 111454
rect 146382 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 217826 111454
rect 218062 111218 218146 111454
rect 218382 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 264250 111454
rect 264486 111218 294970 111454
rect 295206 111218 325690 111454
rect 325926 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 592650 111454
rect -8726 111134 592650 111218
rect -8726 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 73826 111134
rect 74062 110898 74146 111134
rect 74382 110898 109826 111134
rect 110062 110898 110146 111134
rect 110382 110898 145826 111134
rect 146062 110898 146146 111134
rect 146382 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 217826 111134
rect 218062 110898 218146 111134
rect 218382 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 264250 111134
rect 264486 110898 294970 111134
rect 295206 110898 325690 111134
rect 325926 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 592650 111134
rect -8726 110866 592650 110898
rect -8726 106954 592650 106986
rect -8726 106718 -8694 106954
rect -8458 106718 -8374 106954
rect -8138 106718 33326 106954
rect 33562 106718 33646 106954
rect 33882 106718 69326 106954
rect 69562 106718 69646 106954
rect 69882 106718 105326 106954
rect 105562 106718 105646 106954
rect 105882 106718 141326 106954
rect 141562 106718 141646 106954
rect 141882 106718 177326 106954
rect 177562 106718 177646 106954
rect 177882 106718 213326 106954
rect 213562 106718 213646 106954
rect 213882 106718 249326 106954
rect 249562 106718 249646 106954
rect 249882 106718 357326 106954
rect 357562 106718 357646 106954
rect 357882 106718 393326 106954
rect 393562 106718 393646 106954
rect 393882 106718 429326 106954
rect 429562 106718 429646 106954
rect 429882 106718 465326 106954
rect 465562 106718 465646 106954
rect 465882 106718 501326 106954
rect 501562 106718 501646 106954
rect 501882 106718 537326 106954
rect 537562 106718 537646 106954
rect 537882 106718 573326 106954
rect 573562 106718 573646 106954
rect 573882 106718 592062 106954
rect 592298 106718 592382 106954
rect 592618 106718 592650 106954
rect -8726 106634 592650 106718
rect -8726 106398 -8694 106634
rect -8458 106398 -8374 106634
rect -8138 106398 33326 106634
rect 33562 106398 33646 106634
rect 33882 106398 69326 106634
rect 69562 106398 69646 106634
rect 69882 106398 105326 106634
rect 105562 106398 105646 106634
rect 105882 106398 141326 106634
rect 141562 106398 141646 106634
rect 141882 106398 177326 106634
rect 177562 106398 177646 106634
rect 177882 106398 213326 106634
rect 213562 106398 213646 106634
rect 213882 106398 249326 106634
rect 249562 106398 249646 106634
rect 249882 106398 357326 106634
rect 357562 106398 357646 106634
rect 357882 106398 393326 106634
rect 393562 106398 393646 106634
rect 393882 106398 429326 106634
rect 429562 106398 429646 106634
rect 429882 106398 465326 106634
rect 465562 106398 465646 106634
rect 465882 106398 501326 106634
rect 501562 106398 501646 106634
rect 501882 106398 537326 106634
rect 537562 106398 537646 106634
rect 537882 106398 573326 106634
rect 573562 106398 573646 106634
rect 573882 106398 592062 106634
rect 592298 106398 592382 106634
rect 592618 106398 592650 106634
rect -8726 106366 592650 106398
rect -8726 102454 592650 102486
rect -8726 102218 -7734 102454
rect -7498 102218 -7414 102454
rect -7178 102218 28826 102454
rect 29062 102218 29146 102454
rect 29382 102218 64826 102454
rect 65062 102218 65146 102454
rect 65382 102218 100826 102454
rect 101062 102218 101146 102454
rect 101382 102218 136826 102454
rect 137062 102218 137146 102454
rect 137382 102218 172826 102454
rect 173062 102218 173146 102454
rect 173382 102218 208826 102454
rect 209062 102218 209146 102454
rect 209382 102218 244826 102454
rect 245062 102218 245146 102454
rect 245382 102218 352826 102454
rect 353062 102218 353146 102454
rect 353382 102218 388826 102454
rect 389062 102218 389146 102454
rect 389382 102218 424826 102454
rect 425062 102218 425146 102454
rect 425382 102218 460826 102454
rect 461062 102218 461146 102454
rect 461382 102218 496826 102454
rect 497062 102218 497146 102454
rect 497382 102218 532826 102454
rect 533062 102218 533146 102454
rect 533382 102218 568826 102454
rect 569062 102218 569146 102454
rect 569382 102218 591102 102454
rect 591338 102218 591422 102454
rect 591658 102218 592650 102454
rect -8726 102134 592650 102218
rect -8726 101898 -7734 102134
rect -7498 101898 -7414 102134
rect -7178 101898 28826 102134
rect 29062 101898 29146 102134
rect 29382 101898 64826 102134
rect 65062 101898 65146 102134
rect 65382 101898 100826 102134
rect 101062 101898 101146 102134
rect 101382 101898 136826 102134
rect 137062 101898 137146 102134
rect 137382 101898 172826 102134
rect 173062 101898 173146 102134
rect 173382 101898 208826 102134
rect 209062 101898 209146 102134
rect 209382 101898 244826 102134
rect 245062 101898 245146 102134
rect 245382 101898 352826 102134
rect 353062 101898 353146 102134
rect 353382 101898 388826 102134
rect 389062 101898 389146 102134
rect 389382 101898 424826 102134
rect 425062 101898 425146 102134
rect 425382 101898 460826 102134
rect 461062 101898 461146 102134
rect 461382 101898 496826 102134
rect 497062 101898 497146 102134
rect 497382 101898 532826 102134
rect 533062 101898 533146 102134
rect 533382 101898 568826 102134
rect 569062 101898 569146 102134
rect 569382 101898 591102 102134
rect 591338 101898 591422 102134
rect 591658 101898 592650 102134
rect -8726 101866 592650 101898
rect -8726 97954 592650 97986
rect -8726 97718 -6774 97954
rect -6538 97718 -6454 97954
rect -6218 97718 24326 97954
rect 24562 97718 24646 97954
rect 24882 97718 60326 97954
rect 60562 97718 60646 97954
rect 60882 97718 96326 97954
rect 96562 97718 96646 97954
rect 96882 97718 132326 97954
rect 132562 97718 132646 97954
rect 132882 97718 168326 97954
rect 168562 97718 168646 97954
rect 168882 97718 204326 97954
rect 204562 97718 204646 97954
rect 204882 97718 240326 97954
rect 240562 97718 240646 97954
rect 240882 97718 276326 97954
rect 276562 97718 276646 97954
rect 276882 97718 312326 97954
rect 312562 97718 312646 97954
rect 312882 97718 348326 97954
rect 348562 97718 348646 97954
rect 348882 97718 384326 97954
rect 384562 97718 384646 97954
rect 384882 97718 420326 97954
rect 420562 97718 420646 97954
rect 420882 97718 456326 97954
rect 456562 97718 456646 97954
rect 456882 97718 492326 97954
rect 492562 97718 492646 97954
rect 492882 97718 528326 97954
rect 528562 97718 528646 97954
rect 528882 97718 564326 97954
rect 564562 97718 564646 97954
rect 564882 97718 590142 97954
rect 590378 97718 590462 97954
rect 590698 97718 592650 97954
rect -8726 97634 592650 97718
rect -8726 97398 -6774 97634
rect -6538 97398 -6454 97634
rect -6218 97398 24326 97634
rect 24562 97398 24646 97634
rect 24882 97398 60326 97634
rect 60562 97398 60646 97634
rect 60882 97398 96326 97634
rect 96562 97398 96646 97634
rect 96882 97398 132326 97634
rect 132562 97398 132646 97634
rect 132882 97398 168326 97634
rect 168562 97398 168646 97634
rect 168882 97398 204326 97634
rect 204562 97398 204646 97634
rect 204882 97398 240326 97634
rect 240562 97398 240646 97634
rect 240882 97398 276326 97634
rect 276562 97398 276646 97634
rect 276882 97398 312326 97634
rect 312562 97398 312646 97634
rect 312882 97398 348326 97634
rect 348562 97398 348646 97634
rect 348882 97398 384326 97634
rect 384562 97398 384646 97634
rect 384882 97398 420326 97634
rect 420562 97398 420646 97634
rect 420882 97398 456326 97634
rect 456562 97398 456646 97634
rect 456882 97398 492326 97634
rect 492562 97398 492646 97634
rect 492882 97398 528326 97634
rect 528562 97398 528646 97634
rect 528882 97398 564326 97634
rect 564562 97398 564646 97634
rect 564882 97398 590142 97634
rect 590378 97398 590462 97634
rect 590698 97398 592650 97634
rect -8726 97366 592650 97398
rect -8726 93454 592650 93486
rect -8726 93218 -5814 93454
rect -5578 93218 -5494 93454
rect -5258 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 91826 93454
rect 92062 93218 92146 93454
rect 92382 93218 127826 93454
rect 128062 93218 128146 93454
rect 128382 93218 163826 93454
rect 164062 93218 164146 93454
rect 164382 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 589182 93454
rect 589418 93218 589502 93454
rect 589738 93218 592650 93454
rect -8726 93134 592650 93218
rect -8726 92898 -5814 93134
rect -5578 92898 -5494 93134
rect -5258 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 91826 93134
rect 92062 92898 92146 93134
rect 92382 92898 127826 93134
rect 128062 92898 128146 93134
rect 128382 92898 163826 93134
rect 164062 92898 164146 93134
rect 164382 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 589182 93134
rect 589418 92898 589502 93134
rect 589738 92898 592650 93134
rect -8726 92866 592650 92898
rect -8726 88954 592650 88986
rect -8726 88718 -4854 88954
rect -4618 88718 -4534 88954
rect -4298 88718 15326 88954
rect 15562 88718 15646 88954
rect 15882 88718 51326 88954
rect 51562 88718 51646 88954
rect 51882 88718 87326 88954
rect 87562 88718 87646 88954
rect 87882 88718 123326 88954
rect 123562 88718 123646 88954
rect 123882 88718 159326 88954
rect 159562 88718 159646 88954
rect 159882 88718 195326 88954
rect 195562 88718 195646 88954
rect 195882 88718 231326 88954
rect 231562 88718 231646 88954
rect 231882 88718 267326 88954
rect 267562 88718 267646 88954
rect 267882 88718 303326 88954
rect 303562 88718 303646 88954
rect 303882 88718 339326 88954
rect 339562 88718 339646 88954
rect 339882 88718 375326 88954
rect 375562 88718 375646 88954
rect 375882 88718 411326 88954
rect 411562 88718 411646 88954
rect 411882 88718 447326 88954
rect 447562 88718 447646 88954
rect 447882 88718 483326 88954
rect 483562 88718 483646 88954
rect 483882 88718 519326 88954
rect 519562 88718 519646 88954
rect 519882 88718 555326 88954
rect 555562 88718 555646 88954
rect 555882 88718 588222 88954
rect 588458 88718 588542 88954
rect 588778 88718 592650 88954
rect -8726 88634 592650 88718
rect -8726 88398 -4854 88634
rect -4618 88398 -4534 88634
rect -4298 88398 15326 88634
rect 15562 88398 15646 88634
rect 15882 88398 51326 88634
rect 51562 88398 51646 88634
rect 51882 88398 87326 88634
rect 87562 88398 87646 88634
rect 87882 88398 123326 88634
rect 123562 88398 123646 88634
rect 123882 88398 159326 88634
rect 159562 88398 159646 88634
rect 159882 88398 195326 88634
rect 195562 88398 195646 88634
rect 195882 88398 231326 88634
rect 231562 88398 231646 88634
rect 231882 88398 267326 88634
rect 267562 88398 267646 88634
rect 267882 88398 303326 88634
rect 303562 88398 303646 88634
rect 303882 88398 339326 88634
rect 339562 88398 339646 88634
rect 339882 88398 375326 88634
rect 375562 88398 375646 88634
rect 375882 88398 411326 88634
rect 411562 88398 411646 88634
rect 411882 88398 447326 88634
rect 447562 88398 447646 88634
rect 447882 88398 483326 88634
rect 483562 88398 483646 88634
rect 483882 88398 519326 88634
rect 519562 88398 519646 88634
rect 519882 88398 555326 88634
rect 555562 88398 555646 88634
rect 555882 88398 588222 88634
rect 588458 88398 588542 88634
rect 588778 88398 592650 88634
rect -8726 88366 592650 88398
rect -8726 84454 592650 84486
rect -8726 84218 -3894 84454
rect -3658 84218 -3574 84454
rect -3338 84218 10826 84454
rect 11062 84218 11146 84454
rect 11382 84218 46826 84454
rect 47062 84218 47146 84454
rect 47382 84218 82826 84454
rect 83062 84218 83146 84454
rect 83382 84218 118826 84454
rect 119062 84218 119146 84454
rect 119382 84218 154826 84454
rect 155062 84218 155146 84454
rect 155382 84218 190826 84454
rect 191062 84218 191146 84454
rect 191382 84218 226826 84454
rect 227062 84218 227146 84454
rect 227382 84218 262826 84454
rect 263062 84218 263146 84454
rect 263382 84218 298826 84454
rect 299062 84218 299146 84454
rect 299382 84218 334826 84454
rect 335062 84218 335146 84454
rect 335382 84218 370826 84454
rect 371062 84218 371146 84454
rect 371382 84218 406826 84454
rect 407062 84218 407146 84454
rect 407382 84218 442826 84454
rect 443062 84218 443146 84454
rect 443382 84218 478826 84454
rect 479062 84218 479146 84454
rect 479382 84218 514826 84454
rect 515062 84218 515146 84454
rect 515382 84218 550826 84454
rect 551062 84218 551146 84454
rect 551382 84218 587262 84454
rect 587498 84218 587582 84454
rect 587818 84218 592650 84454
rect -8726 84134 592650 84218
rect -8726 83898 -3894 84134
rect -3658 83898 -3574 84134
rect -3338 83898 10826 84134
rect 11062 83898 11146 84134
rect 11382 83898 46826 84134
rect 47062 83898 47146 84134
rect 47382 83898 82826 84134
rect 83062 83898 83146 84134
rect 83382 83898 118826 84134
rect 119062 83898 119146 84134
rect 119382 83898 154826 84134
rect 155062 83898 155146 84134
rect 155382 83898 190826 84134
rect 191062 83898 191146 84134
rect 191382 83898 226826 84134
rect 227062 83898 227146 84134
rect 227382 83898 262826 84134
rect 263062 83898 263146 84134
rect 263382 83898 298826 84134
rect 299062 83898 299146 84134
rect 299382 83898 334826 84134
rect 335062 83898 335146 84134
rect 335382 83898 370826 84134
rect 371062 83898 371146 84134
rect 371382 83898 406826 84134
rect 407062 83898 407146 84134
rect 407382 83898 442826 84134
rect 443062 83898 443146 84134
rect 443382 83898 478826 84134
rect 479062 83898 479146 84134
rect 479382 83898 514826 84134
rect 515062 83898 515146 84134
rect 515382 83898 550826 84134
rect 551062 83898 551146 84134
rect 551382 83898 587262 84134
rect 587498 83898 587582 84134
rect 587818 83898 592650 84134
rect -8726 83866 592650 83898
rect -8726 79954 592650 79986
rect -8726 79718 -2934 79954
rect -2698 79718 -2614 79954
rect -2378 79718 6326 79954
rect 6562 79718 6646 79954
rect 6882 79718 42326 79954
rect 42562 79718 42646 79954
rect 42882 79718 78326 79954
rect 78562 79718 78646 79954
rect 78882 79718 114326 79954
rect 114562 79718 114646 79954
rect 114882 79718 150326 79954
rect 150562 79718 150646 79954
rect 150882 79718 186326 79954
rect 186562 79718 186646 79954
rect 186882 79718 222326 79954
rect 222562 79718 222646 79954
rect 222882 79718 258326 79954
rect 258562 79718 258646 79954
rect 258882 79718 294326 79954
rect 294562 79718 294646 79954
rect 294882 79718 330326 79954
rect 330562 79718 330646 79954
rect 330882 79718 366326 79954
rect 366562 79718 366646 79954
rect 366882 79718 402326 79954
rect 402562 79718 402646 79954
rect 402882 79718 438326 79954
rect 438562 79718 438646 79954
rect 438882 79718 474326 79954
rect 474562 79718 474646 79954
rect 474882 79718 510326 79954
rect 510562 79718 510646 79954
rect 510882 79718 546326 79954
rect 546562 79718 546646 79954
rect 546882 79718 582326 79954
rect 582562 79718 582646 79954
rect 582882 79718 586302 79954
rect 586538 79718 586622 79954
rect 586858 79718 592650 79954
rect -8726 79634 592650 79718
rect -8726 79398 -2934 79634
rect -2698 79398 -2614 79634
rect -2378 79398 6326 79634
rect 6562 79398 6646 79634
rect 6882 79398 42326 79634
rect 42562 79398 42646 79634
rect 42882 79398 78326 79634
rect 78562 79398 78646 79634
rect 78882 79398 114326 79634
rect 114562 79398 114646 79634
rect 114882 79398 150326 79634
rect 150562 79398 150646 79634
rect 150882 79398 186326 79634
rect 186562 79398 186646 79634
rect 186882 79398 222326 79634
rect 222562 79398 222646 79634
rect 222882 79398 258326 79634
rect 258562 79398 258646 79634
rect 258882 79398 294326 79634
rect 294562 79398 294646 79634
rect 294882 79398 330326 79634
rect 330562 79398 330646 79634
rect 330882 79398 366326 79634
rect 366562 79398 366646 79634
rect 366882 79398 402326 79634
rect 402562 79398 402646 79634
rect 402882 79398 438326 79634
rect 438562 79398 438646 79634
rect 438882 79398 474326 79634
rect 474562 79398 474646 79634
rect 474882 79398 510326 79634
rect 510562 79398 510646 79634
rect 510882 79398 546326 79634
rect 546562 79398 546646 79634
rect 546882 79398 582326 79634
rect 582562 79398 582646 79634
rect 582882 79398 586302 79634
rect 586538 79398 586622 79634
rect 586858 79398 592650 79634
rect -8726 79366 592650 79398
rect -8726 75454 592650 75486
rect -8726 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 592650 75454
rect -8726 75134 592650 75218
rect -8726 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 592650 75134
rect -8726 74866 592650 74898
rect -8726 70954 592650 70986
rect -8726 70718 -8694 70954
rect -8458 70718 -8374 70954
rect -8138 70718 33326 70954
rect 33562 70718 33646 70954
rect 33882 70718 69326 70954
rect 69562 70718 69646 70954
rect 69882 70718 105326 70954
rect 105562 70718 105646 70954
rect 105882 70718 141326 70954
rect 141562 70718 141646 70954
rect 141882 70718 177326 70954
rect 177562 70718 177646 70954
rect 177882 70718 213326 70954
rect 213562 70718 213646 70954
rect 213882 70718 249326 70954
rect 249562 70718 249646 70954
rect 249882 70718 285326 70954
rect 285562 70718 285646 70954
rect 285882 70718 321326 70954
rect 321562 70718 321646 70954
rect 321882 70718 357326 70954
rect 357562 70718 357646 70954
rect 357882 70718 393326 70954
rect 393562 70718 393646 70954
rect 393882 70718 429326 70954
rect 429562 70718 429646 70954
rect 429882 70718 465326 70954
rect 465562 70718 465646 70954
rect 465882 70718 501326 70954
rect 501562 70718 501646 70954
rect 501882 70718 537326 70954
rect 537562 70718 537646 70954
rect 537882 70718 573326 70954
rect 573562 70718 573646 70954
rect 573882 70718 592062 70954
rect 592298 70718 592382 70954
rect 592618 70718 592650 70954
rect -8726 70634 592650 70718
rect -8726 70398 -8694 70634
rect -8458 70398 -8374 70634
rect -8138 70398 33326 70634
rect 33562 70398 33646 70634
rect 33882 70398 69326 70634
rect 69562 70398 69646 70634
rect 69882 70398 105326 70634
rect 105562 70398 105646 70634
rect 105882 70398 141326 70634
rect 141562 70398 141646 70634
rect 141882 70398 177326 70634
rect 177562 70398 177646 70634
rect 177882 70398 213326 70634
rect 213562 70398 213646 70634
rect 213882 70398 249326 70634
rect 249562 70398 249646 70634
rect 249882 70398 285326 70634
rect 285562 70398 285646 70634
rect 285882 70398 321326 70634
rect 321562 70398 321646 70634
rect 321882 70398 357326 70634
rect 357562 70398 357646 70634
rect 357882 70398 393326 70634
rect 393562 70398 393646 70634
rect 393882 70398 429326 70634
rect 429562 70398 429646 70634
rect 429882 70398 465326 70634
rect 465562 70398 465646 70634
rect 465882 70398 501326 70634
rect 501562 70398 501646 70634
rect 501882 70398 537326 70634
rect 537562 70398 537646 70634
rect 537882 70398 573326 70634
rect 573562 70398 573646 70634
rect 573882 70398 592062 70634
rect 592298 70398 592382 70634
rect 592618 70398 592650 70634
rect -8726 70366 592650 70398
rect -8726 66454 592650 66486
rect -8726 66218 -7734 66454
rect -7498 66218 -7414 66454
rect -7178 66218 28826 66454
rect 29062 66218 29146 66454
rect 29382 66218 64826 66454
rect 65062 66218 65146 66454
rect 65382 66218 100826 66454
rect 101062 66218 101146 66454
rect 101382 66218 136826 66454
rect 137062 66218 137146 66454
rect 137382 66218 172826 66454
rect 173062 66218 173146 66454
rect 173382 66218 208826 66454
rect 209062 66218 209146 66454
rect 209382 66218 244826 66454
rect 245062 66218 245146 66454
rect 245382 66218 280826 66454
rect 281062 66218 281146 66454
rect 281382 66218 316826 66454
rect 317062 66218 317146 66454
rect 317382 66218 352826 66454
rect 353062 66218 353146 66454
rect 353382 66218 388826 66454
rect 389062 66218 389146 66454
rect 389382 66218 424826 66454
rect 425062 66218 425146 66454
rect 425382 66218 460826 66454
rect 461062 66218 461146 66454
rect 461382 66218 496826 66454
rect 497062 66218 497146 66454
rect 497382 66218 532826 66454
rect 533062 66218 533146 66454
rect 533382 66218 568826 66454
rect 569062 66218 569146 66454
rect 569382 66218 591102 66454
rect 591338 66218 591422 66454
rect 591658 66218 592650 66454
rect -8726 66134 592650 66218
rect -8726 65898 -7734 66134
rect -7498 65898 -7414 66134
rect -7178 65898 28826 66134
rect 29062 65898 29146 66134
rect 29382 65898 64826 66134
rect 65062 65898 65146 66134
rect 65382 65898 100826 66134
rect 101062 65898 101146 66134
rect 101382 65898 136826 66134
rect 137062 65898 137146 66134
rect 137382 65898 172826 66134
rect 173062 65898 173146 66134
rect 173382 65898 208826 66134
rect 209062 65898 209146 66134
rect 209382 65898 244826 66134
rect 245062 65898 245146 66134
rect 245382 65898 280826 66134
rect 281062 65898 281146 66134
rect 281382 65898 316826 66134
rect 317062 65898 317146 66134
rect 317382 65898 352826 66134
rect 353062 65898 353146 66134
rect 353382 65898 388826 66134
rect 389062 65898 389146 66134
rect 389382 65898 424826 66134
rect 425062 65898 425146 66134
rect 425382 65898 460826 66134
rect 461062 65898 461146 66134
rect 461382 65898 496826 66134
rect 497062 65898 497146 66134
rect 497382 65898 532826 66134
rect 533062 65898 533146 66134
rect 533382 65898 568826 66134
rect 569062 65898 569146 66134
rect 569382 65898 591102 66134
rect 591338 65898 591422 66134
rect 591658 65898 592650 66134
rect -8726 65866 592650 65898
rect -8726 61954 592650 61986
rect -8726 61718 -6774 61954
rect -6538 61718 -6454 61954
rect -6218 61718 24326 61954
rect 24562 61718 24646 61954
rect 24882 61718 60326 61954
rect 60562 61718 60646 61954
rect 60882 61718 96326 61954
rect 96562 61718 96646 61954
rect 96882 61718 132326 61954
rect 132562 61718 132646 61954
rect 132882 61718 168326 61954
rect 168562 61718 168646 61954
rect 168882 61718 204326 61954
rect 204562 61718 204646 61954
rect 204882 61718 240326 61954
rect 240562 61718 240646 61954
rect 240882 61718 276326 61954
rect 276562 61718 276646 61954
rect 276882 61718 312326 61954
rect 312562 61718 312646 61954
rect 312882 61718 348326 61954
rect 348562 61718 348646 61954
rect 348882 61718 384326 61954
rect 384562 61718 384646 61954
rect 384882 61718 420326 61954
rect 420562 61718 420646 61954
rect 420882 61718 456326 61954
rect 456562 61718 456646 61954
rect 456882 61718 492326 61954
rect 492562 61718 492646 61954
rect 492882 61718 528326 61954
rect 528562 61718 528646 61954
rect 528882 61718 564326 61954
rect 564562 61718 564646 61954
rect 564882 61718 590142 61954
rect 590378 61718 590462 61954
rect 590698 61718 592650 61954
rect -8726 61634 592650 61718
rect -8726 61398 -6774 61634
rect -6538 61398 -6454 61634
rect -6218 61398 24326 61634
rect 24562 61398 24646 61634
rect 24882 61398 60326 61634
rect 60562 61398 60646 61634
rect 60882 61398 96326 61634
rect 96562 61398 96646 61634
rect 96882 61398 132326 61634
rect 132562 61398 132646 61634
rect 132882 61398 168326 61634
rect 168562 61398 168646 61634
rect 168882 61398 204326 61634
rect 204562 61398 204646 61634
rect 204882 61398 240326 61634
rect 240562 61398 240646 61634
rect 240882 61398 276326 61634
rect 276562 61398 276646 61634
rect 276882 61398 312326 61634
rect 312562 61398 312646 61634
rect 312882 61398 348326 61634
rect 348562 61398 348646 61634
rect 348882 61398 384326 61634
rect 384562 61398 384646 61634
rect 384882 61398 420326 61634
rect 420562 61398 420646 61634
rect 420882 61398 456326 61634
rect 456562 61398 456646 61634
rect 456882 61398 492326 61634
rect 492562 61398 492646 61634
rect 492882 61398 528326 61634
rect 528562 61398 528646 61634
rect 528882 61398 564326 61634
rect 564562 61398 564646 61634
rect 564882 61398 590142 61634
rect 590378 61398 590462 61634
rect 590698 61398 592650 61634
rect -8726 61366 592650 61398
rect -8726 57454 592650 57486
rect -8726 57218 -5814 57454
rect -5578 57218 -5494 57454
rect -5258 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 589182 57454
rect 589418 57218 589502 57454
rect 589738 57218 592650 57454
rect -8726 57134 592650 57218
rect -8726 56898 -5814 57134
rect -5578 56898 -5494 57134
rect -5258 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 589182 57134
rect 589418 56898 589502 57134
rect 589738 56898 592650 57134
rect -8726 56866 592650 56898
rect -8726 52954 592650 52986
rect -8726 52718 -4854 52954
rect -4618 52718 -4534 52954
rect -4298 52718 15326 52954
rect 15562 52718 15646 52954
rect 15882 52718 51326 52954
rect 51562 52718 51646 52954
rect 51882 52718 87326 52954
rect 87562 52718 87646 52954
rect 87882 52718 123326 52954
rect 123562 52718 123646 52954
rect 123882 52718 159326 52954
rect 159562 52718 159646 52954
rect 159882 52718 195326 52954
rect 195562 52718 195646 52954
rect 195882 52718 231326 52954
rect 231562 52718 231646 52954
rect 231882 52718 267326 52954
rect 267562 52718 267646 52954
rect 267882 52718 303326 52954
rect 303562 52718 303646 52954
rect 303882 52718 339326 52954
rect 339562 52718 339646 52954
rect 339882 52718 375326 52954
rect 375562 52718 375646 52954
rect 375882 52718 411326 52954
rect 411562 52718 411646 52954
rect 411882 52718 447326 52954
rect 447562 52718 447646 52954
rect 447882 52718 483326 52954
rect 483562 52718 483646 52954
rect 483882 52718 519326 52954
rect 519562 52718 519646 52954
rect 519882 52718 555326 52954
rect 555562 52718 555646 52954
rect 555882 52718 588222 52954
rect 588458 52718 588542 52954
rect 588778 52718 592650 52954
rect -8726 52634 592650 52718
rect -8726 52398 -4854 52634
rect -4618 52398 -4534 52634
rect -4298 52398 15326 52634
rect 15562 52398 15646 52634
rect 15882 52398 51326 52634
rect 51562 52398 51646 52634
rect 51882 52398 87326 52634
rect 87562 52398 87646 52634
rect 87882 52398 123326 52634
rect 123562 52398 123646 52634
rect 123882 52398 159326 52634
rect 159562 52398 159646 52634
rect 159882 52398 195326 52634
rect 195562 52398 195646 52634
rect 195882 52398 231326 52634
rect 231562 52398 231646 52634
rect 231882 52398 267326 52634
rect 267562 52398 267646 52634
rect 267882 52398 303326 52634
rect 303562 52398 303646 52634
rect 303882 52398 339326 52634
rect 339562 52398 339646 52634
rect 339882 52398 375326 52634
rect 375562 52398 375646 52634
rect 375882 52398 411326 52634
rect 411562 52398 411646 52634
rect 411882 52398 447326 52634
rect 447562 52398 447646 52634
rect 447882 52398 483326 52634
rect 483562 52398 483646 52634
rect 483882 52398 519326 52634
rect 519562 52398 519646 52634
rect 519882 52398 555326 52634
rect 555562 52398 555646 52634
rect 555882 52398 588222 52634
rect 588458 52398 588542 52634
rect 588778 52398 592650 52634
rect -8726 52366 592650 52398
rect -8726 48454 592650 48486
rect -8726 48218 -3894 48454
rect -3658 48218 -3574 48454
rect -3338 48218 10826 48454
rect 11062 48218 11146 48454
rect 11382 48218 46826 48454
rect 47062 48218 47146 48454
rect 47382 48218 82826 48454
rect 83062 48218 83146 48454
rect 83382 48218 118826 48454
rect 119062 48218 119146 48454
rect 119382 48218 154826 48454
rect 155062 48218 155146 48454
rect 155382 48218 190826 48454
rect 191062 48218 191146 48454
rect 191382 48218 226826 48454
rect 227062 48218 227146 48454
rect 227382 48218 262826 48454
rect 263062 48218 263146 48454
rect 263382 48218 298826 48454
rect 299062 48218 299146 48454
rect 299382 48218 334826 48454
rect 335062 48218 335146 48454
rect 335382 48218 370826 48454
rect 371062 48218 371146 48454
rect 371382 48218 406826 48454
rect 407062 48218 407146 48454
rect 407382 48218 442826 48454
rect 443062 48218 443146 48454
rect 443382 48218 478826 48454
rect 479062 48218 479146 48454
rect 479382 48218 514826 48454
rect 515062 48218 515146 48454
rect 515382 48218 550826 48454
rect 551062 48218 551146 48454
rect 551382 48218 587262 48454
rect 587498 48218 587582 48454
rect 587818 48218 592650 48454
rect -8726 48134 592650 48218
rect -8726 47898 -3894 48134
rect -3658 47898 -3574 48134
rect -3338 47898 10826 48134
rect 11062 47898 11146 48134
rect 11382 47898 46826 48134
rect 47062 47898 47146 48134
rect 47382 47898 82826 48134
rect 83062 47898 83146 48134
rect 83382 47898 118826 48134
rect 119062 47898 119146 48134
rect 119382 47898 154826 48134
rect 155062 47898 155146 48134
rect 155382 47898 190826 48134
rect 191062 47898 191146 48134
rect 191382 47898 226826 48134
rect 227062 47898 227146 48134
rect 227382 47898 262826 48134
rect 263062 47898 263146 48134
rect 263382 47898 298826 48134
rect 299062 47898 299146 48134
rect 299382 47898 334826 48134
rect 335062 47898 335146 48134
rect 335382 47898 370826 48134
rect 371062 47898 371146 48134
rect 371382 47898 406826 48134
rect 407062 47898 407146 48134
rect 407382 47898 442826 48134
rect 443062 47898 443146 48134
rect 443382 47898 478826 48134
rect 479062 47898 479146 48134
rect 479382 47898 514826 48134
rect 515062 47898 515146 48134
rect 515382 47898 550826 48134
rect 551062 47898 551146 48134
rect 551382 47898 587262 48134
rect 587498 47898 587582 48134
rect 587818 47898 592650 48134
rect -8726 47866 592650 47898
rect -8726 43954 592650 43986
rect -8726 43718 -2934 43954
rect -2698 43718 -2614 43954
rect -2378 43718 6326 43954
rect 6562 43718 6646 43954
rect 6882 43718 42326 43954
rect 42562 43718 42646 43954
rect 42882 43718 78326 43954
rect 78562 43718 78646 43954
rect 78882 43718 114326 43954
rect 114562 43718 114646 43954
rect 114882 43718 150326 43954
rect 150562 43718 150646 43954
rect 150882 43718 186326 43954
rect 186562 43718 186646 43954
rect 186882 43718 222326 43954
rect 222562 43718 222646 43954
rect 222882 43718 258326 43954
rect 258562 43718 258646 43954
rect 258882 43718 294326 43954
rect 294562 43718 294646 43954
rect 294882 43718 330326 43954
rect 330562 43718 330646 43954
rect 330882 43718 366326 43954
rect 366562 43718 366646 43954
rect 366882 43718 402326 43954
rect 402562 43718 402646 43954
rect 402882 43718 438326 43954
rect 438562 43718 438646 43954
rect 438882 43718 474326 43954
rect 474562 43718 474646 43954
rect 474882 43718 510326 43954
rect 510562 43718 510646 43954
rect 510882 43718 546326 43954
rect 546562 43718 546646 43954
rect 546882 43718 582326 43954
rect 582562 43718 582646 43954
rect 582882 43718 586302 43954
rect 586538 43718 586622 43954
rect 586858 43718 592650 43954
rect -8726 43634 592650 43718
rect -8726 43398 -2934 43634
rect -2698 43398 -2614 43634
rect -2378 43398 6326 43634
rect 6562 43398 6646 43634
rect 6882 43398 42326 43634
rect 42562 43398 42646 43634
rect 42882 43398 78326 43634
rect 78562 43398 78646 43634
rect 78882 43398 114326 43634
rect 114562 43398 114646 43634
rect 114882 43398 150326 43634
rect 150562 43398 150646 43634
rect 150882 43398 186326 43634
rect 186562 43398 186646 43634
rect 186882 43398 222326 43634
rect 222562 43398 222646 43634
rect 222882 43398 258326 43634
rect 258562 43398 258646 43634
rect 258882 43398 294326 43634
rect 294562 43398 294646 43634
rect 294882 43398 330326 43634
rect 330562 43398 330646 43634
rect 330882 43398 366326 43634
rect 366562 43398 366646 43634
rect 366882 43398 402326 43634
rect 402562 43398 402646 43634
rect 402882 43398 438326 43634
rect 438562 43398 438646 43634
rect 438882 43398 474326 43634
rect 474562 43398 474646 43634
rect 474882 43398 510326 43634
rect 510562 43398 510646 43634
rect 510882 43398 546326 43634
rect 546562 43398 546646 43634
rect 546882 43398 582326 43634
rect 582562 43398 582646 43634
rect 582882 43398 586302 43634
rect 586538 43398 586622 43634
rect 586858 43398 592650 43634
rect -8726 43366 592650 43398
rect -8726 39454 592650 39486
rect -8726 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 592650 39454
rect -8726 39134 592650 39218
rect -8726 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 592650 39134
rect -8726 38866 592650 38898
rect -8726 34954 592650 34986
rect -8726 34718 -8694 34954
rect -8458 34718 -8374 34954
rect -8138 34718 33326 34954
rect 33562 34718 33646 34954
rect 33882 34718 69326 34954
rect 69562 34718 69646 34954
rect 69882 34718 105326 34954
rect 105562 34718 105646 34954
rect 105882 34718 141326 34954
rect 141562 34718 141646 34954
rect 141882 34718 177326 34954
rect 177562 34718 177646 34954
rect 177882 34718 213326 34954
rect 213562 34718 213646 34954
rect 213882 34718 249326 34954
rect 249562 34718 249646 34954
rect 249882 34718 285326 34954
rect 285562 34718 285646 34954
rect 285882 34718 321326 34954
rect 321562 34718 321646 34954
rect 321882 34718 357326 34954
rect 357562 34718 357646 34954
rect 357882 34718 393326 34954
rect 393562 34718 393646 34954
rect 393882 34718 429326 34954
rect 429562 34718 429646 34954
rect 429882 34718 465326 34954
rect 465562 34718 465646 34954
rect 465882 34718 501326 34954
rect 501562 34718 501646 34954
rect 501882 34718 537326 34954
rect 537562 34718 537646 34954
rect 537882 34718 573326 34954
rect 573562 34718 573646 34954
rect 573882 34718 592062 34954
rect 592298 34718 592382 34954
rect 592618 34718 592650 34954
rect -8726 34634 592650 34718
rect -8726 34398 -8694 34634
rect -8458 34398 -8374 34634
rect -8138 34398 33326 34634
rect 33562 34398 33646 34634
rect 33882 34398 69326 34634
rect 69562 34398 69646 34634
rect 69882 34398 105326 34634
rect 105562 34398 105646 34634
rect 105882 34398 141326 34634
rect 141562 34398 141646 34634
rect 141882 34398 177326 34634
rect 177562 34398 177646 34634
rect 177882 34398 213326 34634
rect 213562 34398 213646 34634
rect 213882 34398 249326 34634
rect 249562 34398 249646 34634
rect 249882 34398 285326 34634
rect 285562 34398 285646 34634
rect 285882 34398 321326 34634
rect 321562 34398 321646 34634
rect 321882 34398 357326 34634
rect 357562 34398 357646 34634
rect 357882 34398 393326 34634
rect 393562 34398 393646 34634
rect 393882 34398 429326 34634
rect 429562 34398 429646 34634
rect 429882 34398 465326 34634
rect 465562 34398 465646 34634
rect 465882 34398 501326 34634
rect 501562 34398 501646 34634
rect 501882 34398 537326 34634
rect 537562 34398 537646 34634
rect 537882 34398 573326 34634
rect 573562 34398 573646 34634
rect 573882 34398 592062 34634
rect 592298 34398 592382 34634
rect 592618 34398 592650 34634
rect -8726 34366 592650 34398
rect -8726 30454 592650 30486
rect -8726 30218 -7734 30454
rect -7498 30218 -7414 30454
rect -7178 30218 28826 30454
rect 29062 30218 29146 30454
rect 29382 30218 64826 30454
rect 65062 30218 65146 30454
rect 65382 30218 100826 30454
rect 101062 30218 101146 30454
rect 101382 30218 136826 30454
rect 137062 30218 137146 30454
rect 137382 30218 172826 30454
rect 173062 30218 173146 30454
rect 173382 30218 208826 30454
rect 209062 30218 209146 30454
rect 209382 30218 244826 30454
rect 245062 30218 245146 30454
rect 245382 30218 280826 30454
rect 281062 30218 281146 30454
rect 281382 30218 316826 30454
rect 317062 30218 317146 30454
rect 317382 30218 352826 30454
rect 353062 30218 353146 30454
rect 353382 30218 388826 30454
rect 389062 30218 389146 30454
rect 389382 30218 424826 30454
rect 425062 30218 425146 30454
rect 425382 30218 460826 30454
rect 461062 30218 461146 30454
rect 461382 30218 496826 30454
rect 497062 30218 497146 30454
rect 497382 30218 532826 30454
rect 533062 30218 533146 30454
rect 533382 30218 568826 30454
rect 569062 30218 569146 30454
rect 569382 30218 591102 30454
rect 591338 30218 591422 30454
rect 591658 30218 592650 30454
rect -8726 30134 592650 30218
rect -8726 29898 -7734 30134
rect -7498 29898 -7414 30134
rect -7178 29898 28826 30134
rect 29062 29898 29146 30134
rect 29382 29898 64826 30134
rect 65062 29898 65146 30134
rect 65382 29898 100826 30134
rect 101062 29898 101146 30134
rect 101382 29898 136826 30134
rect 137062 29898 137146 30134
rect 137382 29898 172826 30134
rect 173062 29898 173146 30134
rect 173382 29898 208826 30134
rect 209062 29898 209146 30134
rect 209382 29898 244826 30134
rect 245062 29898 245146 30134
rect 245382 29898 280826 30134
rect 281062 29898 281146 30134
rect 281382 29898 316826 30134
rect 317062 29898 317146 30134
rect 317382 29898 352826 30134
rect 353062 29898 353146 30134
rect 353382 29898 388826 30134
rect 389062 29898 389146 30134
rect 389382 29898 424826 30134
rect 425062 29898 425146 30134
rect 425382 29898 460826 30134
rect 461062 29898 461146 30134
rect 461382 29898 496826 30134
rect 497062 29898 497146 30134
rect 497382 29898 532826 30134
rect 533062 29898 533146 30134
rect 533382 29898 568826 30134
rect 569062 29898 569146 30134
rect 569382 29898 591102 30134
rect 591338 29898 591422 30134
rect 591658 29898 592650 30134
rect -8726 29866 592650 29898
rect -8726 25954 592650 25986
rect -8726 25718 -6774 25954
rect -6538 25718 -6454 25954
rect -6218 25718 24326 25954
rect 24562 25718 24646 25954
rect 24882 25718 60326 25954
rect 60562 25718 60646 25954
rect 60882 25718 96326 25954
rect 96562 25718 96646 25954
rect 96882 25718 132326 25954
rect 132562 25718 132646 25954
rect 132882 25718 168326 25954
rect 168562 25718 168646 25954
rect 168882 25718 204326 25954
rect 204562 25718 204646 25954
rect 204882 25718 240326 25954
rect 240562 25718 240646 25954
rect 240882 25718 276326 25954
rect 276562 25718 276646 25954
rect 276882 25718 312326 25954
rect 312562 25718 312646 25954
rect 312882 25718 348326 25954
rect 348562 25718 348646 25954
rect 348882 25718 384326 25954
rect 384562 25718 384646 25954
rect 384882 25718 420326 25954
rect 420562 25718 420646 25954
rect 420882 25718 456326 25954
rect 456562 25718 456646 25954
rect 456882 25718 492326 25954
rect 492562 25718 492646 25954
rect 492882 25718 528326 25954
rect 528562 25718 528646 25954
rect 528882 25718 564326 25954
rect 564562 25718 564646 25954
rect 564882 25718 590142 25954
rect 590378 25718 590462 25954
rect 590698 25718 592650 25954
rect -8726 25634 592650 25718
rect -8726 25398 -6774 25634
rect -6538 25398 -6454 25634
rect -6218 25398 24326 25634
rect 24562 25398 24646 25634
rect 24882 25398 60326 25634
rect 60562 25398 60646 25634
rect 60882 25398 96326 25634
rect 96562 25398 96646 25634
rect 96882 25398 132326 25634
rect 132562 25398 132646 25634
rect 132882 25398 168326 25634
rect 168562 25398 168646 25634
rect 168882 25398 204326 25634
rect 204562 25398 204646 25634
rect 204882 25398 240326 25634
rect 240562 25398 240646 25634
rect 240882 25398 276326 25634
rect 276562 25398 276646 25634
rect 276882 25398 312326 25634
rect 312562 25398 312646 25634
rect 312882 25398 348326 25634
rect 348562 25398 348646 25634
rect 348882 25398 384326 25634
rect 384562 25398 384646 25634
rect 384882 25398 420326 25634
rect 420562 25398 420646 25634
rect 420882 25398 456326 25634
rect 456562 25398 456646 25634
rect 456882 25398 492326 25634
rect 492562 25398 492646 25634
rect 492882 25398 528326 25634
rect 528562 25398 528646 25634
rect 528882 25398 564326 25634
rect 564562 25398 564646 25634
rect 564882 25398 590142 25634
rect 590378 25398 590462 25634
rect 590698 25398 592650 25634
rect -8726 25366 592650 25398
rect -8726 21454 592650 21486
rect -8726 21218 -5814 21454
rect -5578 21218 -5494 21454
rect -5258 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 589182 21454
rect 589418 21218 589502 21454
rect 589738 21218 592650 21454
rect -8726 21134 592650 21218
rect -8726 20898 -5814 21134
rect -5578 20898 -5494 21134
rect -5258 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 589182 21134
rect 589418 20898 589502 21134
rect 589738 20898 592650 21134
rect -8726 20866 592650 20898
rect -8726 16954 592650 16986
rect -8726 16718 -4854 16954
rect -4618 16718 -4534 16954
rect -4298 16718 15326 16954
rect 15562 16718 15646 16954
rect 15882 16718 51326 16954
rect 51562 16718 51646 16954
rect 51882 16718 87326 16954
rect 87562 16718 87646 16954
rect 87882 16718 123326 16954
rect 123562 16718 123646 16954
rect 123882 16718 159326 16954
rect 159562 16718 159646 16954
rect 159882 16718 195326 16954
rect 195562 16718 195646 16954
rect 195882 16718 231326 16954
rect 231562 16718 231646 16954
rect 231882 16718 267326 16954
rect 267562 16718 267646 16954
rect 267882 16718 303326 16954
rect 303562 16718 303646 16954
rect 303882 16718 339326 16954
rect 339562 16718 339646 16954
rect 339882 16718 375326 16954
rect 375562 16718 375646 16954
rect 375882 16718 411326 16954
rect 411562 16718 411646 16954
rect 411882 16718 447326 16954
rect 447562 16718 447646 16954
rect 447882 16718 483326 16954
rect 483562 16718 483646 16954
rect 483882 16718 519326 16954
rect 519562 16718 519646 16954
rect 519882 16718 555326 16954
rect 555562 16718 555646 16954
rect 555882 16718 588222 16954
rect 588458 16718 588542 16954
rect 588778 16718 592650 16954
rect -8726 16634 592650 16718
rect -8726 16398 -4854 16634
rect -4618 16398 -4534 16634
rect -4298 16398 15326 16634
rect 15562 16398 15646 16634
rect 15882 16398 51326 16634
rect 51562 16398 51646 16634
rect 51882 16398 87326 16634
rect 87562 16398 87646 16634
rect 87882 16398 123326 16634
rect 123562 16398 123646 16634
rect 123882 16398 159326 16634
rect 159562 16398 159646 16634
rect 159882 16398 195326 16634
rect 195562 16398 195646 16634
rect 195882 16398 231326 16634
rect 231562 16398 231646 16634
rect 231882 16398 267326 16634
rect 267562 16398 267646 16634
rect 267882 16398 303326 16634
rect 303562 16398 303646 16634
rect 303882 16398 339326 16634
rect 339562 16398 339646 16634
rect 339882 16398 375326 16634
rect 375562 16398 375646 16634
rect 375882 16398 411326 16634
rect 411562 16398 411646 16634
rect 411882 16398 447326 16634
rect 447562 16398 447646 16634
rect 447882 16398 483326 16634
rect 483562 16398 483646 16634
rect 483882 16398 519326 16634
rect 519562 16398 519646 16634
rect 519882 16398 555326 16634
rect 555562 16398 555646 16634
rect 555882 16398 588222 16634
rect 588458 16398 588542 16634
rect 588778 16398 592650 16634
rect -8726 16366 592650 16398
rect -8726 12454 592650 12486
rect -8726 12218 -3894 12454
rect -3658 12218 -3574 12454
rect -3338 12218 10826 12454
rect 11062 12218 11146 12454
rect 11382 12218 46826 12454
rect 47062 12218 47146 12454
rect 47382 12218 82826 12454
rect 83062 12218 83146 12454
rect 83382 12218 118826 12454
rect 119062 12218 119146 12454
rect 119382 12218 154826 12454
rect 155062 12218 155146 12454
rect 155382 12218 190826 12454
rect 191062 12218 191146 12454
rect 191382 12218 226826 12454
rect 227062 12218 227146 12454
rect 227382 12218 262826 12454
rect 263062 12218 263146 12454
rect 263382 12218 298826 12454
rect 299062 12218 299146 12454
rect 299382 12218 334826 12454
rect 335062 12218 335146 12454
rect 335382 12218 370826 12454
rect 371062 12218 371146 12454
rect 371382 12218 406826 12454
rect 407062 12218 407146 12454
rect 407382 12218 442826 12454
rect 443062 12218 443146 12454
rect 443382 12218 478826 12454
rect 479062 12218 479146 12454
rect 479382 12218 514826 12454
rect 515062 12218 515146 12454
rect 515382 12218 550826 12454
rect 551062 12218 551146 12454
rect 551382 12218 587262 12454
rect 587498 12218 587582 12454
rect 587818 12218 592650 12454
rect -8726 12134 592650 12218
rect -8726 11898 -3894 12134
rect -3658 11898 -3574 12134
rect -3338 11898 10826 12134
rect 11062 11898 11146 12134
rect 11382 11898 46826 12134
rect 47062 11898 47146 12134
rect 47382 11898 82826 12134
rect 83062 11898 83146 12134
rect 83382 11898 118826 12134
rect 119062 11898 119146 12134
rect 119382 11898 154826 12134
rect 155062 11898 155146 12134
rect 155382 11898 190826 12134
rect 191062 11898 191146 12134
rect 191382 11898 226826 12134
rect 227062 11898 227146 12134
rect 227382 11898 262826 12134
rect 263062 11898 263146 12134
rect 263382 11898 298826 12134
rect 299062 11898 299146 12134
rect 299382 11898 334826 12134
rect 335062 11898 335146 12134
rect 335382 11898 370826 12134
rect 371062 11898 371146 12134
rect 371382 11898 406826 12134
rect 407062 11898 407146 12134
rect 407382 11898 442826 12134
rect 443062 11898 443146 12134
rect 443382 11898 478826 12134
rect 479062 11898 479146 12134
rect 479382 11898 514826 12134
rect 515062 11898 515146 12134
rect 515382 11898 550826 12134
rect 551062 11898 551146 12134
rect 551382 11898 587262 12134
rect 587498 11898 587582 12134
rect 587818 11898 592650 12134
rect -8726 11866 592650 11898
rect -8726 7954 592650 7986
rect -8726 7718 -2934 7954
rect -2698 7718 -2614 7954
rect -2378 7718 6326 7954
rect 6562 7718 6646 7954
rect 6882 7718 42326 7954
rect 42562 7718 42646 7954
rect 42882 7718 78326 7954
rect 78562 7718 78646 7954
rect 78882 7718 114326 7954
rect 114562 7718 114646 7954
rect 114882 7718 150326 7954
rect 150562 7718 150646 7954
rect 150882 7718 186326 7954
rect 186562 7718 186646 7954
rect 186882 7718 222326 7954
rect 222562 7718 222646 7954
rect 222882 7718 258326 7954
rect 258562 7718 258646 7954
rect 258882 7718 294326 7954
rect 294562 7718 294646 7954
rect 294882 7718 330326 7954
rect 330562 7718 330646 7954
rect 330882 7718 366326 7954
rect 366562 7718 366646 7954
rect 366882 7718 402326 7954
rect 402562 7718 402646 7954
rect 402882 7718 438326 7954
rect 438562 7718 438646 7954
rect 438882 7718 474326 7954
rect 474562 7718 474646 7954
rect 474882 7718 510326 7954
rect 510562 7718 510646 7954
rect 510882 7718 546326 7954
rect 546562 7718 546646 7954
rect 546882 7718 582326 7954
rect 582562 7718 582646 7954
rect 582882 7718 586302 7954
rect 586538 7718 586622 7954
rect 586858 7718 592650 7954
rect -8726 7634 592650 7718
rect -8726 7398 -2934 7634
rect -2698 7398 -2614 7634
rect -2378 7398 6326 7634
rect 6562 7398 6646 7634
rect 6882 7398 42326 7634
rect 42562 7398 42646 7634
rect 42882 7398 78326 7634
rect 78562 7398 78646 7634
rect 78882 7398 114326 7634
rect 114562 7398 114646 7634
rect 114882 7398 150326 7634
rect 150562 7398 150646 7634
rect 150882 7398 186326 7634
rect 186562 7398 186646 7634
rect 186882 7398 222326 7634
rect 222562 7398 222646 7634
rect 222882 7398 258326 7634
rect 258562 7398 258646 7634
rect 258882 7398 294326 7634
rect 294562 7398 294646 7634
rect 294882 7398 330326 7634
rect 330562 7398 330646 7634
rect 330882 7398 366326 7634
rect 366562 7398 366646 7634
rect 366882 7398 402326 7634
rect 402562 7398 402646 7634
rect 402882 7398 438326 7634
rect 438562 7398 438646 7634
rect 438882 7398 474326 7634
rect 474562 7398 474646 7634
rect 474882 7398 510326 7634
rect 510562 7398 510646 7634
rect 510882 7398 546326 7634
rect 546562 7398 546646 7634
rect 546882 7398 582326 7634
rect 582562 7398 582646 7634
rect 582882 7398 586302 7634
rect 586538 7398 586622 7634
rect 586858 7398 592650 7634
rect -8726 7366 592650 7398
rect -8726 3454 592650 3486
rect -8726 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 592650 3454
rect -8726 3134 592650 3218
rect -8726 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 592650 3134
rect -8726 2866 592650 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 6326 -1306
rect 6562 -1542 6646 -1306
rect 6882 -1542 42326 -1306
rect 42562 -1542 42646 -1306
rect 42882 -1542 78326 -1306
rect 78562 -1542 78646 -1306
rect 78882 -1542 114326 -1306
rect 114562 -1542 114646 -1306
rect 114882 -1542 150326 -1306
rect 150562 -1542 150646 -1306
rect 150882 -1542 186326 -1306
rect 186562 -1542 186646 -1306
rect 186882 -1542 222326 -1306
rect 222562 -1542 222646 -1306
rect 222882 -1542 258326 -1306
rect 258562 -1542 258646 -1306
rect 258882 -1542 294326 -1306
rect 294562 -1542 294646 -1306
rect 294882 -1542 330326 -1306
rect 330562 -1542 330646 -1306
rect 330882 -1542 366326 -1306
rect 366562 -1542 366646 -1306
rect 366882 -1542 402326 -1306
rect 402562 -1542 402646 -1306
rect 402882 -1542 438326 -1306
rect 438562 -1542 438646 -1306
rect 438882 -1542 474326 -1306
rect 474562 -1542 474646 -1306
rect 474882 -1542 510326 -1306
rect 510562 -1542 510646 -1306
rect 510882 -1542 546326 -1306
rect 546562 -1542 546646 -1306
rect 546882 -1542 582326 -1306
rect 582562 -1542 582646 -1306
rect 582882 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 6326 -1626
rect 6562 -1862 6646 -1626
rect 6882 -1862 42326 -1626
rect 42562 -1862 42646 -1626
rect 42882 -1862 78326 -1626
rect 78562 -1862 78646 -1626
rect 78882 -1862 114326 -1626
rect 114562 -1862 114646 -1626
rect 114882 -1862 150326 -1626
rect 150562 -1862 150646 -1626
rect 150882 -1862 186326 -1626
rect 186562 -1862 186646 -1626
rect 186882 -1862 222326 -1626
rect 222562 -1862 222646 -1626
rect 222882 -1862 258326 -1626
rect 258562 -1862 258646 -1626
rect 258882 -1862 294326 -1626
rect 294562 -1862 294646 -1626
rect 294882 -1862 330326 -1626
rect 330562 -1862 330646 -1626
rect 330882 -1862 366326 -1626
rect 366562 -1862 366646 -1626
rect 366882 -1862 402326 -1626
rect 402562 -1862 402646 -1626
rect 402882 -1862 438326 -1626
rect 438562 -1862 438646 -1626
rect 438882 -1862 474326 -1626
rect 474562 -1862 474646 -1626
rect 474882 -1862 510326 -1626
rect 510562 -1862 510646 -1626
rect 510882 -1862 546326 -1626
rect 546562 -1862 546646 -1626
rect 546882 -1862 582326 -1626
rect 582562 -1862 582646 -1626
rect 582882 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 10826 -2266
rect 11062 -2502 11146 -2266
rect 11382 -2502 46826 -2266
rect 47062 -2502 47146 -2266
rect 47382 -2502 82826 -2266
rect 83062 -2502 83146 -2266
rect 83382 -2502 118826 -2266
rect 119062 -2502 119146 -2266
rect 119382 -2502 154826 -2266
rect 155062 -2502 155146 -2266
rect 155382 -2502 190826 -2266
rect 191062 -2502 191146 -2266
rect 191382 -2502 226826 -2266
rect 227062 -2502 227146 -2266
rect 227382 -2502 262826 -2266
rect 263062 -2502 263146 -2266
rect 263382 -2502 298826 -2266
rect 299062 -2502 299146 -2266
rect 299382 -2502 334826 -2266
rect 335062 -2502 335146 -2266
rect 335382 -2502 370826 -2266
rect 371062 -2502 371146 -2266
rect 371382 -2502 406826 -2266
rect 407062 -2502 407146 -2266
rect 407382 -2502 442826 -2266
rect 443062 -2502 443146 -2266
rect 443382 -2502 478826 -2266
rect 479062 -2502 479146 -2266
rect 479382 -2502 514826 -2266
rect 515062 -2502 515146 -2266
rect 515382 -2502 550826 -2266
rect 551062 -2502 551146 -2266
rect 551382 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 10826 -2586
rect 11062 -2822 11146 -2586
rect 11382 -2822 46826 -2586
rect 47062 -2822 47146 -2586
rect 47382 -2822 82826 -2586
rect 83062 -2822 83146 -2586
rect 83382 -2822 118826 -2586
rect 119062 -2822 119146 -2586
rect 119382 -2822 154826 -2586
rect 155062 -2822 155146 -2586
rect 155382 -2822 190826 -2586
rect 191062 -2822 191146 -2586
rect 191382 -2822 226826 -2586
rect 227062 -2822 227146 -2586
rect 227382 -2822 262826 -2586
rect 263062 -2822 263146 -2586
rect 263382 -2822 298826 -2586
rect 299062 -2822 299146 -2586
rect 299382 -2822 334826 -2586
rect 335062 -2822 335146 -2586
rect 335382 -2822 370826 -2586
rect 371062 -2822 371146 -2586
rect 371382 -2822 406826 -2586
rect 407062 -2822 407146 -2586
rect 407382 -2822 442826 -2586
rect 443062 -2822 443146 -2586
rect 443382 -2822 478826 -2586
rect 479062 -2822 479146 -2586
rect 479382 -2822 514826 -2586
rect 515062 -2822 515146 -2586
rect 515382 -2822 550826 -2586
rect 551062 -2822 551146 -2586
rect 551382 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 15326 -3226
rect 15562 -3462 15646 -3226
rect 15882 -3462 51326 -3226
rect 51562 -3462 51646 -3226
rect 51882 -3462 87326 -3226
rect 87562 -3462 87646 -3226
rect 87882 -3462 123326 -3226
rect 123562 -3462 123646 -3226
rect 123882 -3462 159326 -3226
rect 159562 -3462 159646 -3226
rect 159882 -3462 195326 -3226
rect 195562 -3462 195646 -3226
rect 195882 -3462 231326 -3226
rect 231562 -3462 231646 -3226
rect 231882 -3462 267326 -3226
rect 267562 -3462 267646 -3226
rect 267882 -3462 303326 -3226
rect 303562 -3462 303646 -3226
rect 303882 -3462 339326 -3226
rect 339562 -3462 339646 -3226
rect 339882 -3462 375326 -3226
rect 375562 -3462 375646 -3226
rect 375882 -3462 411326 -3226
rect 411562 -3462 411646 -3226
rect 411882 -3462 447326 -3226
rect 447562 -3462 447646 -3226
rect 447882 -3462 483326 -3226
rect 483562 -3462 483646 -3226
rect 483882 -3462 519326 -3226
rect 519562 -3462 519646 -3226
rect 519882 -3462 555326 -3226
rect 555562 -3462 555646 -3226
rect 555882 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 15326 -3546
rect 15562 -3782 15646 -3546
rect 15882 -3782 51326 -3546
rect 51562 -3782 51646 -3546
rect 51882 -3782 87326 -3546
rect 87562 -3782 87646 -3546
rect 87882 -3782 123326 -3546
rect 123562 -3782 123646 -3546
rect 123882 -3782 159326 -3546
rect 159562 -3782 159646 -3546
rect 159882 -3782 195326 -3546
rect 195562 -3782 195646 -3546
rect 195882 -3782 231326 -3546
rect 231562 -3782 231646 -3546
rect 231882 -3782 267326 -3546
rect 267562 -3782 267646 -3546
rect 267882 -3782 303326 -3546
rect 303562 -3782 303646 -3546
rect 303882 -3782 339326 -3546
rect 339562 -3782 339646 -3546
rect 339882 -3782 375326 -3546
rect 375562 -3782 375646 -3546
rect 375882 -3782 411326 -3546
rect 411562 -3782 411646 -3546
rect 411882 -3782 447326 -3546
rect 447562 -3782 447646 -3546
rect 447882 -3782 483326 -3546
rect 483562 -3782 483646 -3546
rect 483882 -3782 519326 -3546
rect 519562 -3782 519646 -3546
rect 519882 -3782 555326 -3546
rect 555562 -3782 555646 -3546
rect 555882 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 19826 -4186
rect 20062 -4422 20146 -4186
rect 20382 -4422 55826 -4186
rect 56062 -4422 56146 -4186
rect 56382 -4422 91826 -4186
rect 92062 -4422 92146 -4186
rect 92382 -4422 127826 -4186
rect 128062 -4422 128146 -4186
rect 128382 -4422 163826 -4186
rect 164062 -4422 164146 -4186
rect 164382 -4422 199826 -4186
rect 200062 -4422 200146 -4186
rect 200382 -4422 235826 -4186
rect 236062 -4422 236146 -4186
rect 236382 -4422 271826 -4186
rect 272062 -4422 272146 -4186
rect 272382 -4422 307826 -4186
rect 308062 -4422 308146 -4186
rect 308382 -4422 343826 -4186
rect 344062 -4422 344146 -4186
rect 344382 -4422 379826 -4186
rect 380062 -4422 380146 -4186
rect 380382 -4422 415826 -4186
rect 416062 -4422 416146 -4186
rect 416382 -4422 451826 -4186
rect 452062 -4422 452146 -4186
rect 452382 -4422 487826 -4186
rect 488062 -4422 488146 -4186
rect 488382 -4422 523826 -4186
rect 524062 -4422 524146 -4186
rect 524382 -4422 559826 -4186
rect 560062 -4422 560146 -4186
rect 560382 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 19826 -4506
rect 20062 -4742 20146 -4506
rect 20382 -4742 55826 -4506
rect 56062 -4742 56146 -4506
rect 56382 -4742 91826 -4506
rect 92062 -4742 92146 -4506
rect 92382 -4742 127826 -4506
rect 128062 -4742 128146 -4506
rect 128382 -4742 163826 -4506
rect 164062 -4742 164146 -4506
rect 164382 -4742 199826 -4506
rect 200062 -4742 200146 -4506
rect 200382 -4742 235826 -4506
rect 236062 -4742 236146 -4506
rect 236382 -4742 271826 -4506
rect 272062 -4742 272146 -4506
rect 272382 -4742 307826 -4506
rect 308062 -4742 308146 -4506
rect 308382 -4742 343826 -4506
rect 344062 -4742 344146 -4506
rect 344382 -4742 379826 -4506
rect 380062 -4742 380146 -4506
rect 380382 -4742 415826 -4506
rect 416062 -4742 416146 -4506
rect 416382 -4742 451826 -4506
rect 452062 -4742 452146 -4506
rect 452382 -4742 487826 -4506
rect 488062 -4742 488146 -4506
rect 488382 -4742 523826 -4506
rect 524062 -4742 524146 -4506
rect 524382 -4742 559826 -4506
rect 560062 -4742 560146 -4506
rect 560382 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 24326 -5146
rect 24562 -5382 24646 -5146
rect 24882 -5382 60326 -5146
rect 60562 -5382 60646 -5146
rect 60882 -5382 96326 -5146
rect 96562 -5382 96646 -5146
rect 96882 -5382 132326 -5146
rect 132562 -5382 132646 -5146
rect 132882 -5382 168326 -5146
rect 168562 -5382 168646 -5146
rect 168882 -5382 204326 -5146
rect 204562 -5382 204646 -5146
rect 204882 -5382 240326 -5146
rect 240562 -5382 240646 -5146
rect 240882 -5382 276326 -5146
rect 276562 -5382 276646 -5146
rect 276882 -5382 312326 -5146
rect 312562 -5382 312646 -5146
rect 312882 -5382 348326 -5146
rect 348562 -5382 348646 -5146
rect 348882 -5382 384326 -5146
rect 384562 -5382 384646 -5146
rect 384882 -5382 420326 -5146
rect 420562 -5382 420646 -5146
rect 420882 -5382 456326 -5146
rect 456562 -5382 456646 -5146
rect 456882 -5382 492326 -5146
rect 492562 -5382 492646 -5146
rect 492882 -5382 528326 -5146
rect 528562 -5382 528646 -5146
rect 528882 -5382 564326 -5146
rect 564562 -5382 564646 -5146
rect 564882 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 24326 -5466
rect 24562 -5702 24646 -5466
rect 24882 -5702 60326 -5466
rect 60562 -5702 60646 -5466
rect 60882 -5702 96326 -5466
rect 96562 -5702 96646 -5466
rect 96882 -5702 132326 -5466
rect 132562 -5702 132646 -5466
rect 132882 -5702 168326 -5466
rect 168562 -5702 168646 -5466
rect 168882 -5702 204326 -5466
rect 204562 -5702 204646 -5466
rect 204882 -5702 240326 -5466
rect 240562 -5702 240646 -5466
rect 240882 -5702 276326 -5466
rect 276562 -5702 276646 -5466
rect 276882 -5702 312326 -5466
rect 312562 -5702 312646 -5466
rect 312882 -5702 348326 -5466
rect 348562 -5702 348646 -5466
rect 348882 -5702 384326 -5466
rect 384562 -5702 384646 -5466
rect 384882 -5702 420326 -5466
rect 420562 -5702 420646 -5466
rect 420882 -5702 456326 -5466
rect 456562 -5702 456646 -5466
rect 456882 -5702 492326 -5466
rect 492562 -5702 492646 -5466
rect 492882 -5702 528326 -5466
rect 528562 -5702 528646 -5466
rect 528882 -5702 564326 -5466
rect 564562 -5702 564646 -5466
rect 564882 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 28826 -6106
rect 29062 -6342 29146 -6106
rect 29382 -6342 64826 -6106
rect 65062 -6342 65146 -6106
rect 65382 -6342 100826 -6106
rect 101062 -6342 101146 -6106
rect 101382 -6342 136826 -6106
rect 137062 -6342 137146 -6106
rect 137382 -6342 172826 -6106
rect 173062 -6342 173146 -6106
rect 173382 -6342 208826 -6106
rect 209062 -6342 209146 -6106
rect 209382 -6342 244826 -6106
rect 245062 -6342 245146 -6106
rect 245382 -6342 280826 -6106
rect 281062 -6342 281146 -6106
rect 281382 -6342 316826 -6106
rect 317062 -6342 317146 -6106
rect 317382 -6342 352826 -6106
rect 353062 -6342 353146 -6106
rect 353382 -6342 388826 -6106
rect 389062 -6342 389146 -6106
rect 389382 -6342 424826 -6106
rect 425062 -6342 425146 -6106
rect 425382 -6342 460826 -6106
rect 461062 -6342 461146 -6106
rect 461382 -6342 496826 -6106
rect 497062 -6342 497146 -6106
rect 497382 -6342 532826 -6106
rect 533062 -6342 533146 -6106
rect 533382 -6342 568826 -6106
rect 569062 -6342 569146 -6106
rect 569382 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 28826 -6426
rect 29062 -6662 29146 -6426
rect 29382 -6662 64826 -6426
rect 65062 -6662 65146 -6426
rect 65382 -6662 100826 -6426
rect 101062 -6662 101146 -6426
rect 101382 -6662 136826 -6426
rect 137062 -6662 137146 -6426
rect 137382 -6662 172826 -6426
rect 173062 -6662 173146 -6426
rect 173382 -6662 208826 -6426
rect 209062 -6662 209146 -6426
rect 209382 -6662 244826 -6426
rect 245062 -6662 245146 -6426
rect 245382 -6662 280826 -6426
rect 281062 -6662 281146 -6426
rect 281382 -6662 316826 -6426
rect 317062 -6662 317146 -6426
rect 317382 -6662 352826 -6426
rect 353062 -6662 353146 -6426
rect 353382 -6662 388826 -6426
rect 389062 -6662 389146 -6426
rect 389382 -6662 424826 -6426
rect 425062 -6662 425146 -6426
rect 425382 -6662 460826 -6426
rect 461062 -6662 461146 -6426
rect 461382 -6662 496826 -6426
rect 497062 -6662 497146 -6426
rect 497382 -6662 532826 -6426
rect 533062 -6662 533146 -6426
rect 533382 -6662 568826 -6426
rect 569062 -6662 569146 -6426
rect 569382 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 33326 -7066
rect 33562 -7302 33646 -7066
rect 33882 -7302 69326 -7066
rect 69562 -7302 69646 -7066
rect 69882 -7302 105326 -7066
rect 105562 -7302 105646 -7066
rect 105882 -7302 141326 -7066
rect 141562 -7302 141646 -7066
rect 141882 -7302 177326 -7066
rect 177562 -7302 177646 -7066
rect 177882 -7302 213326 -7066
rect 213562 -7302 213646 -7066
rect 213882 -7302 249326 -7066
rect 249562 -7302 249646 -7066
rect 249882 -7302 285326 -7066
rect 285562 -7302 285646 -7066
rect 285882 -7302 321326 -7066
rect 321562 -7302 321646 -7066
rect 321882 -7302 357326 -7066
rect 357562 -7302 357646 -7066
rect 357882 -7302 393326 -7066
rect 393562 -7302 393646 -7066
rect 393882 -7302 429326 -7066
rect 429562 -7302 429646 -7066
rect 429882 -7302 465326 -7066
rect 465562 -7302 465646 -7066
rect 465882 -7302 501326 -7066
rect 501562 -7302 501646 -7066
rect 501882 -7302 537326 -7066
rect 537562 -7302 537646 -7066
rect 537882 -7302 573326 -7066
rect 573562 -7302 573646 -7066
rect 573882 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 33326 -7386
rect 33562 -7622 33646 -7386
rect 33882 -7622 69326 -7386
rect 69562 -7622 69646 -7386
rect 69882 -7622 105326 -7386
rect 105562 -7622 105646 -7386
rect 105882 -7622 141326 -7386
rect 141562 -7622 141646 -7386
rect 141882 -7622 177326 -7386
rect 177562 -7622 177646 -7386
rect 177882 -7622 213326 -7386
rect 213562 -7622 213646 -7386
rect 213882 -7622 249326 -7386
rect 249562 -7622 249646 -7386
rect 249882 -7622 285326 -7386
rect 285562 -7622 285646 -7386
rect 285882 -7622 321326 -7386
rect 321562 -7622 321646 -7386
rect 321882 -7622 357326 -7386
rect 357562 -7622 357646 -7386
rect 357882 -7622 393326 -7386
rect 393562 -7622 393646 -7386
rect 393882 -7622 429326 -7386
rect 429562 -7622 429646 -7386
rect 429882 -7622 465326 -7386
rect 465562 -7622 465646 -7386
rect 465882 -7622 501326 -7386
rect 501562 -7622 501646 -7386
rect 501882 -7622 537326 -7386
rect 537562 -7622 537646 -7386
rect 537882 -7622 573326 -7386
rect 573562 -7622 573646 -7386
rect 573882 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use cpu  cpu0
timestamp 0
transform 1 0 260000 0 1 100000
box 0 0 84000 56000
use sky130_sram_1kbyte_1rw1r_8x1024_8  memHword
timestamp 0
transform 1 0 380000 0 1 500000
box 0 0 91060 89292
use sky130_sram_1kbyte_1rw1r_8x1024_8  memLword
timestamp 0
transform 1 0 100000 0 1 500000
box 0 0 91060 89292
use soc_config  mprj
timestamp 0
transform 1 0 235000 0 1 338000
box 1066 0 64898 44000
<< labels >>
flabel metal3 s 583520 285276 584960 285516 0 FreeSans 960 0 0 0 analog_io[0]
port 0 nsew signal bidirectional
flabel metal2 s 446098 703520 446210 704960 0 FreeSans 448 90 0 0 analog_io[10]
port 1 nsew signal bidirectional
flabel metal2 s 381146 703520 381258 704960 0 FreeSans 448 90 0 0 analog_io[11]
port 2 nsew signal bidirectional
flabel metal2 s 316286 703520 316398 704960 0 FreeSans 448 90 0 0 analog_io[12]
port 3 nsew signal bidirectional
flabel metal2 s 251426 703520 251538 704960 0 FreeSans 448 90 0 0 analog_io[13]
port 4 nsew signal bidirectional
flabel metal2 s 186474 703520 186586 704960 0 FreeSans 448 90 0 0 analog_io[14]
port 5 nsew signal bidirectional
flabel metal2 s 121614 703520 121726 704960 0 FreeSans 448 90 0 0 analog_io[15]
port 6 nsew signal bidirectional
flabel metal2 s 56754 703520 56866 704960 0 FreeSans 448 90 0 0 analog_io[16]
port 7 nsew signal bidirectional
flabel metal3 s -960 697220 480 697460 0 FreeSans 960 0 0 0 analog_io[17]
port 8 nsew signal bidirectional
flabel metal3 s -960 644996 480 645236 0 FreeSans 960 0 0 0 analog_io[18]
port 9 nsew signal bidirectional
flabel metal3 s -960 592908 480 593148 0 FreeSans 960 0 0 0 analog_io[19]
port 10 nsew signal bidirectional
flabel metal3 s 583520 338452 584960 338692 0 FreeSans 960 0 0 0 analog_io[1]
port 11 nsew signal bidirectional
flabel metal3 s -960 540684 480 540924 0 FreeSans 960 0 0 0 analog_io[20]
port 12 nsew signal bidirectional
flabel metal3 s -960 488596 480 488836 0 FreeSans 960 0 0 0 analog_io[21]
port 13 nsew signal bidirectional
flabel metal3 s -960 436508 480 436748 0 FreeSans 960 0 0 0 analog_io[22]
port 14 nsew signal bidirectional
flabel metal3 s -960 384284 480 384524 0 FreeSans 960 0 0 0 analog_io[23]
port 15 nsew signal bidirectional
flabel metal3 s -960 332196 480 332436 0 FreeSans 960 0 0 0 analog_io[24]
port 16 nsew signal bidirectional
flabel metal3 s -960 279972 480 280212 0 FreeSans 960 0 0 0 analog_io[25]
port 17 nsew signal bidirectional
flabel metal3 s -960 227884 480 228124 0 FreeSans 960 0 0 0 analog_io[26]
port 18 nsew signal bidirectional
flabel metal3 s -960 175796 480 176036 0 FreeSans 960 0 0 0 analog_io[27]
port 19 nsew signal bidirectional
flabel metal3 s -960 123572 480 123812 0 FreeSans 960 0 0 0 analog_io[28]
port 20 nsew signal bidirectional
flabel metal3 s 583520 391628 584960 391868 0 FreeSans 960 0 0 0 analog_io[2]
port 21 nsew signal bidirectional
flabel metal3 s 583520 444668 584960 444908 0 FreeSans 960 0 0 0 analog_io[3]
port 22 nsew signal bidirectional
flabel metal3 s 583520 497844 584960 498084 0 FreeSans 960 0 0 0 analog_io[4]
port 23 nsew signal bidirectional
flabel metal3 s 583520 551020 584960 551260 0 FreeSans 960 0 0 0 analog_io[5]
port 24 nsew signal bidirectional
flabel metal3 s 583520 604060 584960 604300 0 FreeSans 960 0 0 0 analog_io[6]
port 25 nsew signal bidirectional
flabel metal3 s 583520 657236 584960 657476 0 FreeSans 960 0 0 0 analog_io[7]
port 26 nsew signal bidirectional
flabel metal2 s 575818 703520 575930 704960 0 FreeSans 448 90 0 0 analog_io[8]
port 27 nsew signal bidirectional
flabel metal2 s 510958 703520 511070 704960 0 FreeSans 448 90 0 0 analog_io[9]
port 28 nsew signal bidirectional
flabel metal3 s 583520 6476 584960 6716 0 FreeSans 960 0 0 0 io_in[0]
port 29 nsew signal input
flabel metal3 s 583520 457996 584960 458236 0 FreeSans 960 0 0 0 io_in[10]
port 30 nsew signal input
flabel metal3 s 583520 511172 584960 511412 0 FreeSans 960 0 0 0 io_in[11]
port 31 nsew signal input
flabel metal3 s 583520 564212 584960 564452 0 FreeSans 960 0 0 0 io_in[12]
port 32 nsew signal input
flabel metal3 s 583520 617388 584960 617628 0 FreeSans 960 0 0 0 io_in[13]
port 33 nsew signal input
flabel metal3 s 583520 670564 584960 670804 0 FreeSans 960 0 0 0 io_in[14]
port 34 nsew signal input
flabel metal2 s 559626 703520 559738 704960 0 FreeSans 448 90 0 0 io_in[15]
port 35 nsew signal input
flabel metal2 s 494766 703520 494878 704960 0 FreeSans 448 90 0 0 io_in[16]
port 36 nsew signal input
flabel metal2 s 429814 703520 429926 704960 0 FreeSans 448 90 0 0 io_in[17]
port 37 nsew signal input
flabel metal2 s 364954 703520 365066 704960 0 FreeSans 448 90 0 0 io_in[18]
port 38 nsew signal input
flabel metal2 s 300094 703520 300206 704960 0 FreeSans 448 90 0 0 io_in[19]
port 39 nsew signal input
flabel metal3 s 583520 46188 584960 46428 0 FreeSans 960 0 0 0 io_in[1]
port 40 nsew signal input
flabel metal2 s 235142 703520 235254 704960 0 FreeSans 448 90 0 0 io_in[20]
port 41 nsew signal input
flabel metal2 s 170282 703520 170394 704960 0 FreeSans 448 90 0 0 io_in[21]
port 42 nsew signal input
flabel metal2 s 105422 703520 105534 704960 0 FreeSans 448 90 0 0 io_in[22]
port 43 nsew signal input
flabel metal2 s 40470 703520 40582 704960 0 FreeSans 448 90 0 0 io_in[23]
port 44 nsew signal input
flabel metal3 s -960 684164 480 684404 0 FreeSans 960 0 0 0 io_in[24]
port 45 nsew signal input
flabel metal3 s -960 631940 480 632180 0 FreeSans 960 0 0 0 io_in[25]
port 46 nsew signal input
flabel metal3 s -960 579852 480 580092 0 FreeSans 960 0 0 0 io_in[26]
port 47 nsew signal input
flabel metal3 s -960 527764 480 528004 0 FreeSans 960 0 0 0 io_in[27]
port 48 nsew signal input
flabel metal3 s -960 475540 480 475780 0 FreeSans 960 0 0 0 io_in[28]
port 49 nsew signal input
flabel metal3 s -960 423452 480 423692 0 FreeSans 960 0 0 0 io_in[29]
port 50 nsew signal input
flabel metal3 s 583520 86036 584960 86276 0 FreeSans 960 0 0 0 io_in[2]
port 51 nsew signal input
flabel metal3 s -960 371228 480 371468 0 FreeSans 960 0 0 0 io_in[30]
port 52 nsew signal input
flabel metal3 s -960 319140 480 319380 0 FreeSans 960 0 0 0 io_in[31]
port 53 nsew signal input
flabel metal3 s -960 267052 480 267292 0 FreeSans 960 0 0 0 io_in[32]
port 54 nsew signal input
flabel metal3 s -960 214828 480 215068 0 FreeSans 960 0 0 0 io_in[33]
port 55 nsew signal input
flabel metal3 s -960 162740 480 162980 0 FreeSans 960 0 0 0 io_in[34]
port 56 nsew signal input
flabel metal3 s -960 110516 480 110756 0 FreeSans 960 0 0 0 io_in[35]
port 57 nsew signal input
flabel metal3 s -960 71484 480 71724 0 FreeSans 960 0 0 0 io_in[36]
port 58 nsew signal input
flabel metal3 s -960 32316 480 32556 0 FreeSans 960 0 0 0 io_in[37]
port 59 nsew signal input
flabel metal3 s 583520 125884 584960 126124 0 FreeSans 960 0 0 0 io_in[3]
port 60 nsew signal input
flabel metal3 s 583520 165732 584960 165972 0 FreeSans 960 0 0 0 io_in[4]
port 61 nsew signal input
flabel metal3 s 583520 205580 584960 205820 0 FreeSans 960 0 0 0 io_in[5]
port 62 nsew signal input
flabel metal3 s 583520 245428 584960 245668 0 FreeSans 960 0 0 0 io_in[6]
port 63 nsew signal input
flabel metal3 s 583520 298604 584960 298844 0 FreeSans 960 0 0 0 io_in[7]
port 64 nsew signal input
flabel metal3 s 583520 351780 584960 352020 0 FreeSans 960 0 0 0 io_in[8]
port 65 nsew signal input
flabel metal3 s 583520 404820 584960 405060 0 FreeSans 960 0 0 0 io_in[9]
port 66 nsew signal input
flabel metal3 s 583520 32996 584960 33236 0 FreeSans 960 0 0 0 io_oeb[0]
port 67 nsew signal tristate
flabel metal3 s 583520 484516 584960 484756 0 FreeSans 960 0 0 0 io_oeb[10]
port 68 nsew signal tristate
flabel metal3 s 583520 537692 584960 537932 0 FreeSans 960 0 0 0 io_oeb[11]
port 69 nsew signal tristate
flabel metal3 s 583520 590868 584960 591108 0 FreeSans 960 0 0 0 io_oeb[12]
port 70 nsew signal tristate
flabel metal3 s 583520 643908 584960 644148 0 FreeSans 960 0 0 0 io_oeb[13]
port 71 nsew signal tristate
flabel metal3 s 583520 697084 584960 697324 0 FreeSans 960 0 0 0 io_oeb[14]
port 72 nsew signal tristate
flabel metal2 s 527150 703520 527262 704960 0 FreeSans 448 90 0 0 io_oeb[15]
port 73 nsew signal tristate
flabel metal2 s 462290 703520 462402 704960 0 FreeSans 448 90 0 0 io_oeb[16]
port 74 nsew signal tristate
flabel metal2 s 397430 703520 397542 704960 0 FreeSans 448 90 0 0 io_oeb[17]
port 75 nsew signal tristate
flabel metal2 s 332478 703520 332590 704960 0 FreeSans 448 90 0 0 io_oeb[18]
port 76 nsew signal tristate
flabel metal2 s 267618 703520 267730 704960 0 FreeSans 448 90 0 0 io_oeb[19]
port 77 nsew signal tristate
flabel metal3 s 583520 72844 584960 73084 0 FreeSans 960 0 0 0 io_oeb[1]
port 78 nsew signal tristate
flabel metal2 s 202758 703520 202870 704960 0 FreeSans 448 90 0 0 io_oeb[20]
port 79 nsew signal tristate
flabel metal2 s 137806 703520 137918 704960 0 FreeSans 448 90 0 0 io_oeb[21]
port 80 nsew signal tristate
flabel metal2 s 72946 703520 73058 704960 0 FreeSans 448 90 0 0 io_oeb[22]
port 81 nsew signal tristate
flabel metal2 s 8086 703520 8198 704960 0 FreeSans 448 90 0 0 io_oeb[23]
port 82 nsew signal tristate
flabel metal3 s -960 658052 480 658292 0 FreeSans 960 0 0 0 io_oeb[24]
port 83 nsew signal tristate
flabel metal3 s -960 605964 480 606204 0 FreeSans 960 0 0 0 io_oeb[25]
port 84 nsew signal tristate
flabel metal3 s -960 553740 480 553980 0 FreeSans 960 0 0 0 io_oeb[26]
port 85 nsew signal tristate
flabel metal3 s -960 501652 480 501892 0 FreeSans 960 0 0 0 io_oeb[27]
port 86 nsew signal tristate
flabel metal3 s -960 449428 480 449668 0 FreeSans 960 0 0 0 io_oeb[28]
port 87 nsew signal tristate
flabel metal3 s -960 397340 480 397580 0 FreeSans 960 0 0 0 io_oeb[29]
port 88 nsew signal tristate
flabel metal3 s 583520 112692 584960 112932 0 FreeSans 960 0 0 0 io_oeb[2]
port 89 nsew signal tristate
flabel metal3 s -960 345252 480 345492 0 FreeSans 960 0 0 0 io_oeb[30]
port 90 nsew signal tristate
flabel metal3 s -960 293028 480 293268 0 FreeSans 960 0 0 0 io_oeb[31]
port 91 nsew signal tristate
flabel metal3 s -960 240940 480 241180 0 FreeSans 960 0 0 0 io_oeb[32]
port 92 nsew signal tristate
flabel metal3 s -960 188716 480 188956 0 FreeSans 960 0 0 0 io_oeb[33]
port 93 nsew signal tristate
flabel metal3 s -960 136628 480 136868 0 FreeSans 960 0 0 0 io_oeb[34]
port 94 nsew signal tristate
flabel metal3 s -960 84540 480 84780 0 FreeSans 960 0 0 0 io_oeb[35]
port 95 nsew signal tristate
flabel metal3 s -960 45372 480 45612 0 FreeSans 960 0 0 0 io_oeb[36]
port 96 nsew signal tristate
flabel metal3 s -960 6340 480 6580 0 FreeSans 960 0 0 0 io_oeb[37]
port 97 nsew signal tristate
flabel metal3 s 583520 152540 584960 152780 0 FreeSans 960 0 0 0 io_oeb[3]
port 98 nsew signal tristate
flabel metal3 s 583520 192388 584960 192628 0 FreeSans 960 0 0 0 io_oeb[4]
port 99 nsew signal tristate
flabel metal3 s 583520 232236 584960 232476 0 FreeSans 960 0 0 0 io_oeb[5]
port 100 nsew signal tristate
flabel metal3 s 583520 272084 584960 272324 0 FreeSans 960 0 0 0 io_oeb[6]
port 101 nsew signal tristate
flabel metal3 s 583520 325124 584960 325364 0 FreeSans 960 0 0 0 io_oeb[7]
port 102 nsew signal tristate
flabel metal3 s 583520 378300 584960 378540 0 FreeSans 960 0 0 0 io_oeb[8]
port 103 nsew signal tristate
flabel metal3 s 583520 431476 584960 431716 0 FreeSans 960 0 0 0 io_oeb[9]
port 104 nsew signal tristate
flabel metal3 s 583520 19668 584960 19908 0 FreeSans 960 0 0 0 io_out[0]
port 105 nsew signal tristate
flabel metal3 s 583520 471324 584960 471564 0 FreeSans 960 0 0 0 io_out[10]
port 106 nsew signal tristate
flabel metal3 s 583520 524364 584960 524604 0 FreeSans 960 0 0 0 io_out[11]
port 107 nsew signal tristate
flabel metal3 s 583520 577540 584960 577780 0 FreeSans 960 0 0 0 io_out[12]
port 108 nsew signal tristate
flabel metal3 s 583520 630716 584960 630956 0 FreeSans 960 0 0 0 io_out[13]
port 109 nsew signal tristate
flabel metal3 s 583520 683756 584960 683996 0 FreeSans 960 0 0 0 io_out[14]
port 110 nsew signal tristate
flabel metal2 s 543434 703520 543546 704960 0 FreeSans 448 90 0 0 io_out[15]
port 111 nsew signal tristate
flabel metal2 s 478482 703520 478594 704960 0 FreeSans 448 90 0 0 io_out[16]
port 112 nsew signal tristate
flabel metal2 s 413622 703520 413734 704960 0 FreeSans 448 90 0 0 io_out[17]
port 113 nsew signal tristate
flabel metal2 s 348762 703520 348874 704960 0 FreeSans 448 90 0 0 io_out[18]
port 114 nsew signal tristate
flabel metal2 s 283810 703520 283922 704960 0 FreeSans 448 90 0 0 io_out[19]
port 115 nsew signal tristate
flabel metal3 s 583520 59516 584960 59756 0 FreeSans 960 0 0 0 io_out[1]
port 116 nsew signal tristate
flabel metal2 s 218950 703520 219062 704960 0 FreeSans 448 90 0 0 io_out[20]
port 117 nsew signal tristate
flabel metal2 s 154090 703520 154202 704960 0 FreeSans 448 90 0 0 io_out[21]
port 118 nsew signal tristate
flabel metal2 s 89138 703520 89250 704960 0 FreeSans 448 90 0 0 io_out[22]
port 119 nsew signal tristate
flabel metal2 s 24278 703520 24390 704960 0 FreeSans 448 90 0 0 io_out[23]
port 120 nsew signal tristate
flabel metal3 s -960 671108 480 671348 0 FreeSans 960 0 0 0 io_out[24]
port 121 nsew signal tristate
flabel metal3 s -960 619020 480 619260 0 FreeSans 960 0 0 0 io_out[25]
port 122 nsew signal tristate
flabel metal3 s -960 566796 480 567036 0 FreeSans 960 0 0 0 io_out[26]
port 123 nsew signal tristate
flabel metal3 s -960 514708 480 514948 0 FreeSans 960 0 0 0 io_out[27]
port 124 nsew signal tristate
flabel metal3 s -960 462484 480 462724 0 FreeSans 960 0 0 0 io_out[28]
port 125 nsew signal tristate
flabel metal3 s -960 410396 480 410636 0 FreeSans 960 0 0 0 io_out[29]
port 126 nsew signal tristate
flabel metal3 s 583520 99364 584960 99604 0 FreeSans 960 0 0 0 io_out[2]
port 127 nsew signal tristate
flabel metal3 s -960 358308 480 358548 0 FreeSans 960 0 0 0 io_out[30]
port 128 nsew signal tristate
flabel metal3 s -960 306084 480 306324 0 FreeSans 960 0 0 0 io_out[31]
port 129 nsew signal tristate
flabel metal3 s -960 253996 480 254236 0 FreeSans 960 0 0 0 io_out[32]
port 130 nsew signal tristate
flabel metal3 s -960 201772 480 202012 0 FreeSans 960 0 0 0 io_out[33]
port 131 nsew signal tristate
flabel metal3 s -960 149684 480 149924 0 FreeSans 960 0 0 0 io_out[34]
port 132 nsew signal tristate
flabel metal3 s -960 97460 480 97700 0 FreeSans 960 0 0 0 io_out[35]
port 133 nsew signal tristate
flabel metal3 s -960 58428 480 58668 0 FreeSans 960 0 0 0 io_out[36]
port 134 nsew signal tristate
flabel metal3 s -960 19260 480 19500 0 FreeSans 960 0 0 0 io_out[37]
port 135 nsew signal tristate
flabel metal3 s 583520 139212 584960 139452 0 FreeSans 960 0 0 0 io_out[3]
port 136 nsew signal tristate
flabel metal3 s 583520 179060 584960 179300 0 FreeSans 960 0 0 0 io_out[4]
port 137 nsew signal tristate
flabel metal3 s 583520 218908 584960 219148 0 FreeSans 960 0 0 0 io_out[5]
port 138 nsew signal tristate
flabel metal3 s 583520 258756 584960 258996 0 FreeSans 960 0 0 0 io_out[6]
port 139 nsew signal tristate
flabel metal3 s 583520 311932 584960 312172 0 FreeSans 960 0 0 0 io_out[7]
port 140 nsew signal tristate
flabel metal3 s 583520 364972 584960 365212 0 FreeSans 960 0 0 0 io_out[8]
port 141 nsew signal tristate
flabel metal3 s 583520 418148 584960 418388 0 FreeSans 960 0 0 0 io_out[9]
port 142 nsew signal tristate
flabel metal2 s 125846 -960 125958 480 0 FreeSans 448 90 0 0 la_data_in[0]
port 143 nsew signal input
flabel metal2 s 480506 -960 480618 480 0 FreeSans 448 90 0 0 la_data_in[100]
port 144 nsew signal input
flabel metal2 s 484002 -960 484114 480 0 FreeSans 448 90 0 0 la_data_in[101]
port 145 nsew signal input
flabel metal2 s 487590 -960 487702 480 0 FreeSans 448 90 0 0 la_data_in[102]
port 146 nsew signal input
flabel metal2 s 491086 -960 491198 480 0 FreeSans 448 90 0 0 la_data_in[103]
port 147 nsew signal input
flabel metal2 s 494674 -960 494786 480 0 FreeSans 448 90 0 0 la_data_in[104]
port 148 nsew signal input
flabel metal2 s 498170 -960 498282 480 0 FreeSans 448 90 0 0 la_data_in[105]
port 149 nsew signal input
flabel metal2 s 501758 -960 501870 480 0 FreeSans 448 90 0 0 la_data_in[106]
port 150 nsew signal input
flabel metal2 s 505346 -960 505458 480 0 FreeSans 448 90 0 0 la_data_in[107]
port 151 nsew signal input
flabel metal2 s 508842 -960 508954 480 0 FreeSans 448 90 0 0 la_data_in[108]
port 152 nsew signal input
flabel metal2 s 512430 -960 512542 480 0 FreeSans 448 90 0 0 la_data_in[109]
port 153 nsew signal input
flabel metal2 s 161266 -960 161378 480 0 FreeSans 448 90 0 0 la_data_in[10]
port 154 nsew signal input
flabel metal2 s 515926 -960 516038 480 0 FreeSans 448 90 0 0 la_data_in[110]
port 155 nsew signal input
flabel metal2 s 519514 -960 519626 480 0 FreeSans 448 90 0 0 la_data_in[111]
port 156 nsew signal input
flabel metal2 s 523010 -960 523122 480 0 FreeSans 448 90 0 0 la_data_in[112]
port 157 nsew signal input
flabel metal2 s 526598 -960 526710 480 0 FreeSans 448 90 0 0 la_data_in[113]
port 158 nsew signal input
flabel metal2 s 530094 -960 530206 480 0 FreeSans 448 90 0 0 la_data_in[114]
port 159 nsew signal input
flabel metal2 s 533682 -960 533794 480 0 FreeSans 448 90 0 0 la_data_in[115]
port 160 nsew signal input
flabel metal2 s 537178 -960 537290 480 0 FreeSans 448 90 0 0 la_data_in[116]
port 161 nsew signal input
flabel metal2 s 540766 -960 540878 480 0 FreeSans 448 90 0 0 la_data_in[117]
port 162 nsew signal input
flabel metal2 s 544354 -960 544466 480 0 FreeSans 448 90 0 0 la_data_in[118]
port 163 nsew signal input
flabel metal2 s 547850 -960 547962 480 0 FreeSans 448 90 0 0 la_data_in[119]
port 164 nsew signal input
flabel metal2 s 164854 -960 164966 480 0 FreeSans 448 90 0 0 la_data_in[11]
port 165 nsew signal input
flabel metal2 s 551438 -960 551550 480 0 FreeSans 448 90 0 0 la_data_in[120]
port 166 nsew signal input
flabel metal2 s 554934 -960 555046 480 0 FreeSans 448 90 0 0 la_data_in[121]
port 167 nsew signal input
flabel metal2 s 558522 -960 558634 480 0 FreeSans 448 90 0 0 la_data_in[122]
port 168 nsew signal input
flabel metal2 s 562018 -960 562130 480 0 FreeSans 448 90 0 0 la_data_in[123]
port 169 nsew signal input
flabel metal2 s 565606 -960 565718 480 0 FreeSans 448 90 0 0 la_data_in[124]
port 170 nsew signal input
flabel metal2 s 569102 -960 569214 480 0 FreeSans 448 90 0 0 la_data_in[125]
port 171 nsew signal input
flabel metal2 s 572690 -960 572802 480 0 FreeSans 448 90 0 0 la_data_in[126]
port 172 nsew signal input
flabel metal2 s 576278 -960 576390 480 0 FreeSans 448 90 0 0 la_data_in[127]
port 173 nsew signal input
flabel metal2 s 168350 -960 168462 480 0 FreeSans 448 90 0 0 la_data_in[12]
port 174 nsew signal input
flabel metal2 s 171938 -960 172050 480 0 FreeSans 448 90 0 0 la_data_in[13]
port 175 nsew signal input
flabel metal2 s 175434 -960 175546 480 0 FreeSans 448 90 0 0 la_data_in[14]
port 176 nsew signal input
flabel metal2 s 179022 -960 179134 480 0 FreeSans 448 90 0 0 la_data_in[15]
port 177 nsew signal input
flabel metal2 s 182518 -960 182630 480 0 FreeSans 448 90 0 0 la_data_in[16]
port 178 nsew signal input
flabel metal2 s 186106 -960 186218 480 0 FreeSans 448 90 0 0 la_data_in[17]
port 179 nsew signal input
flabel metal2 s 189694 -960 189806 480 0 FreeSans 448 90 0 0 la_data_in[18]
port 180 nsew signal input
flabel metal2 s 193190 -960 193302 480 0 FreeSans 448 90 0 0 la_data_in[19]
port 181 nsew signal input
flabel metal2 s 129342 -960 129454 480 0 FreeSans 448 90 0 0 la_data_in[1]
port 182 nsew signal input
flabel metal2 s 196778 -960 196890 480 0 FreeSans 448 90 0 0 la_data_in[20]
port 183 nsew signal input
flabel metal2 s 200274 -960 200386 480 0 FreeSans 448 90 0 0 la_data_in[21]
port 184 nsew signal input
flabel metal2 s 203862 -960 203974 480 0 FreeSans 448 90 0 0 la_data_in[22]
port 185 nsew signal input
flabel metal2 s 207358 -960 207470 480 0 FreeSans 448 90 0 0 la_data_in[23]
port 186 nsew signal input
flabel metal2 s 210946 -960 211058 480 0 FreeSans 448 90 0 0 la_data_in[24]
port 187 nsew signal input
flabel metal2 s 214442 -960 214554 480 0 FreeSans 448 90 0 0 la_data_in[25]
port 188 nsew signal input
flabel metal2 s 218030 -960 218142 480 0 FreeSans 448 90 0 0 la_data_in[26]
port 189 nsew signal input
flabel metal2 s 221526 -960 221638 480 0 FreeSans 448 90 0 0 la_data_in[27]
port 190 nsew signal input
flabel metal2 s 225114 -960 225226 480 0 FreeSans 448 90 0 0 la_data_in[28]
port 191 nsew signal input
flabel metal2 s 228702 -960 228814 480 0 FreeSans 448 90 0 0 la_data_in[29]
port 192 nsew signal input
flabel metal2 s 132930 -960 133042 480 0 FreeSans 448 90 0 0 la_data_in[2]
port 193 nsew signal input
flabel metal2 s 232198 -960 232310 480 0 FreeSans 448 90 0 0 la_data_in[30]
port 194 nsew signal input
flabel metal2 s 235786 -960 235898 480 0 FreeSans 448 90 0 0 la_data_in[31]
port 195 nsew signal input
flabel metal2 s 239282 -960 239394 480 0 FreeSans 448 90 0 0 la_data_in[32]
port 196 nsew signal input
flabel metal2 s 242870 -960 242982 480 0 FreeSans 448 90 0 0 la_data_in[33]
port 197 nsew signal input
flabel metal2 s 246366 -960 246478 480 0 FreeSans 448 90 0 0 la_data_in[34]
port 198 nsew signal input
flabel metal2 s 249954 -960 250066 480 0 FreeSans 448 90 0 0 la_data_in[35]
port 199 nsew signal input
flabel metal2 s 253450 -960 253562 480 0 FreeSans 448 90 0 0 la_data_in[36]
port 200 nsew signal input
flabel metal2 s 257038 -960 257150 480 0 FreeSans 448 90 0 0 la_data_in[37]
port 201 nsew signal input
flabel metal2 s 260626 -960 260738 480 0 FreeSans 448 90 0 0 la_data_in[38]
port 202 nsew signal input
flabel metal2 s 264122 -960 264234 480 0 FreeSans 448 90 0 0 la_data_in[39]
port 203 nsew signal input
flabel metal2 s 136426 -960 136538 480 0 FreeSans 448 90 0 0 la_data_in[3]
port 204 nsew signal input
flabel metal2 s 267710 -960 267822 480 0 FreeSans 448 90 0 0 la_data_in[40]
port 205 nsew signal input
flabel metal2 s 271206 -960 271318 480 0 FreeSans 448 90 0 0 la_data_in[41]
port 206 nsew signal input
flabel metal2 s 274794 -960 274906 480 0 FreeSans 448 90 0 0 la_data_in[42]
port 207 nsew signal input
flabel metal2 s 278290 -960 278402 480 0 FreeSans 448 90 0 0 la_data_in[43]
port 208 nsew signal input
flabel metal2 s 281878 -960 281990 480 0 FreeSans 448 90 0 0 la_data_in[44]
port 209 nsew signal input
flabel metal2 s 285374 -960 285486 480 0 FreeSans 448 90 0 0 la_data_in[45]
port 210 nsew signal input
flabel metal2 s 288962 -960 289074 480 0 FreeSans 448 90 0 0 la_data_in[46]
port 211 nsew signal input
flabel metal2 s 292550 -960 292662 480 0 FreeSans 448 90 0 0 la_data_in[47]
port 212 nsew signal input
flabel metal2 s 296046 -960 296158 480 0 FreeSans 448 90 0 0 la_data_in[48]
port 213 nsew signal input
flabel metal2 s 299634 -960 299746 480 0 FreeSans 448 90 0 0 la_data_in[49]
port 214 nsew signal input
flabel metal2 s 140014 -960 140126 480 0 FreeSans 448 90 0 0 la_data_in[4]
port 215 nsew signal input
flabel metal2 s 303130 -960 303242 480 0 FreeSans 448 90 0 0 la_data_in[50]
port 216 nsew signal input
flabel metal2 s 306718 -960 306830 480 0 FreeSans 448 90 0 0 la_data_in[51]
port 217 nsew signal input
flabel metal2 s 310214 -960 310326 480 0 FreeSans 448 90 0 0 la_data_in[52]
port 218 nsew signal input
flabel metal2 s 313802 -960 313914 480 0 FreeSans 448 90 0 0 la_data_in[53]
port 219 nsew signal input
flabel metal2 s 317298 -960 317410 480 0 FreeSans 448 90 0 0 la_data_in[54]
port 220 nsew signal input
flabel metal2 s 320886 -960 320998 480 0 FreeSans 448 90 0 0 la_data_in[55]
port 221 nsew signal input
flabel metal2 s 324382 -960 324494 480 0 FreeSans 448 90 0 0 la_data_in[56]
port 222 nsew signal input
flabel metal2 s 327970 -960 328082 480 0 FreeSans 448 90 0 0 la_data_in[57]
port 223 nsew signal input
flabel metal2 s 331558 -960 331670 480 0 FreeSans 448 90 0 0 la_data_in[58]
port 224 nsew signal input
flabel metal2 s 335054 -960 335166 480 0 FreeSans 448 90 0 0 la_data_in[59]
port 225 nsew signal input
flabel metal2 s 143510 -960 143622 480 0 FreeSans 448 90 0 0 la_data_in[5]
port 226 nsew signal input
flabel metal2 s 338642 -960 338754 480 0 FreeSans 448 90 0 0 la_data_in[60]
port 227 nsew signal input
flabel metal2 s 342138 -960 342250 480 0 FreeSans 448 90 0 0 la_data_in[61]
port 228 nsew signal input
flabel metal2 s 345726 -960 345838 480 0 FreeSans 448 90 0 0 la_data_in[62]
port 229 nsew signal input
flabel metal2 s 349222 -960 349334 480 0 FreeSans 448 90 0 0 la_data_in[63]
port 230 nsew signal input
flabel metal2 s 352810 -960 352922 480 0 FreeSans 448 90 0 0 la_data_in[64]
port 231 nsew signal input
flabel metal2 s 356306 -960 356418 480 0 FreeSans 448 90 0 0 la_data_in[65]
port 232 nsew signal input
flabel metal2 s 359894 -960 360006 480 0 FreeSans 448 90 0 0 la_data_in[66]
port 233 nsew signal input
flabel metal2 s 363482 -960 363594 480 0 FreeSans 448 90 0 0 la_data_in[67]
port 234 nsew signal input
flabel metal2 s 366978 -960 367090 480 0 FreeSans 448 90 0 0 la_data_in[68]
port 235 nsew signal input
flabel metal2 s 370566 -960 370678 480 0 FreeSans 448 90 0 0 la_data_in[69]
port 236 nsew signal input
flabel metal2 s 147098 -960 147210 480 0 FreeSans 448 90 0 0 la_data_in[6]
port 237 nsew signal input
flabel metal2 s 374062 -960 374174 480 0 FreeSans 448 90 0 0 la_data_in[70]
port 238 nsew signal input
flabel metal2 s 377650 -960 377762 480 0 FreeSans 448 90 0 0 la_data_in[71]
port 239 nsew signal input
flabel metal2 s 381146 -960 381258 480 0 FreeSans 448 90 0 0 la_data_in[72]
port 240 nsew signal input
flabel metal2 s 384734 -960 384846 480 0 FreeSans 448 90 0 0 la_data_in[73]
port 241 nsew signal input
flabel metal2 s 388230 -960 388342 480 0 FreeSans 448 90 0 0 la_data_in[74]
port 242 nsew signal input
flabel metal2 s 391818 -960 391930 480 0 FreeSans 448 90 0 0 la_data_in[75]
port 243 nsew signal input
flabel metal2 s 395314 -960 395426 480 0 FreeSans 448 90 0 0 la_data_in[76]
port 244 nsew signal input
flabel metal2 s 398902 -960 399014 480 0 FreeSans 448 90 0 0 la_data_in[77]
port 245 nsew signal input
flabel metal2 s 402490 -960 402602 480 0 FreeSans 448 90 0 0 la_data_in[78]
port 246 nsew signal input
flabel metal2 s 405986 -960 406098 480 0 FreeSans 448 90 0 0 la_data_in[79]
port 247 nsew signal input
flabel metal2 s 150594 -960 150706 480 0 FreeSans 448 90 0 0 la_data_in[7]
port 248 nsew signal input
flabel metal2 s 409574 -960 409686 480 0 FreeSans 448 90 0 0 la_data_in[80]
port 249 nsew signal input
flabel metal2 s 413070 -960 413182 480 0 FreeSans 448 90 0 0 la_data_in[81]
port 250 nsew signal input
flabel metal2 s 416658 -960 416770 480 0 FreeSans 448 90 0 0 la_data_in[82]
port 251 nsew signal input
flabel metal2 s 420154 -960 420266 480 0 FreeSans 448 90 0 0 la_data_in[83]
port 252 nsew signal input
flabel metal2 s 423742 -960 423854 480 0 FreeSans 448 90 0 0 la_data_in[84]
port 253 nsew signal input
flabel metal2 s 427238 -960 427350 480 0 FreeSans 448 90 0 0 la_data_in[85]
port 254 nsew signal input
flabel metal2 s 430826 -960 430938 480 0 FreeSans 448 90 0 0 la_data_in[86]
port 255 nsew signal input
flabel metal2 s 434414 -960 434526 480 0 FreeSans 448 90 0 0 la_data_in[87]
port 256 nsew signal input
flabel metal2 s 437910 -960 438022 480 0 FreeSans 448 90 0 0 la_data_in[88]
port 257 nsew signal input
flabel metal2 s 441498 -960 441610 480 0 FreeSans 448 90 0 0 la_data_in[89]
port 258 nsew signal input
flabel metal2 s 154182 -960 154294 480 0 FreeSans 448 90 0 0 la_data_in[8]
port 259 nsew signal input
flabel metal2 s 444994 -960 445106 480 0 FreeSans 448 90 0 0 la_data_in[90]
port 260 nsew signal input
flabel metal2 s 448582 -960 448694 480 0 FreeSans 448 90 0 0 la_data_in[91]
port 261 nsew signal input
flabel metal2 s 452078 -960 452190 480 0 FreeSans 448 90 0 0 la_data_in[92]
port 262 nsew signal input
flabel metal2 s 455666 -960 455778 480 0 FreeSans 448 90 0 0 la_data_in[93]
port 263 nsew signal input
flabel metal2 s 459162 -960 459274 480 0 FreeSans 448 90 0 0 la_data_in[94]
port 264 nsew signal input
flabel metal2 s 462750 -960 462862 480 0 FreeSans 448 90 0 0 la_data_in[95]
port 265 nsew signal input
flabel metal2 s 466246 -960 466358 480 0 FreeSans 448 90 0 0 la_data_in[96]
port 266 nsew signal input
flabel metal2 s 469834 -960 469946 480 0 FreeSans 448 90 0 0 la_data_in[97]
port 267 nsew signal input
flabel metal2 s 473422 -960 473534 480 0 FreeSans 448 90 0 0 la_data_in[98]
port 268 nsew signal input
flabel metal2 s 476918 -960 477030 480 0 FreeSans 448 90 0 0 la_data_in[99]
port 269 nsew signal input
flabel metal2 s 157770 -960 157882 480 0 FreeSans 448 90 0 0 la_data_in[9]
port 270 nsew signal input
flabel metal2 s 126950 -960 127062 480 0 FreeSans 448 90 0 0 la_data_out[0]
port 271 nsew signal tristate
flabel metal2 s 481702 -960 481814 480 0 FreeSans 448 90 0 0 la_data_out[100]
port 272 nsew signal tristate
flabel metal2 s 485198 -960 485310 480 0 FreeSans 448 90 0 0 la_data_out[101]
port 273 nsew signal tristate
flabel metal2 s 488786 -960 488898 480 0 FreeSans 448 90 0 0 la_data_out[102]
port 274 nsew signal tristate
flabel metal2 s 492282 -960 492394 480 0 FreeSans 448 90 0 0 la_data_out[103]
port 275 nsew signal tristate
flabel metal2 s 495870 -960 495982 480 0 FreeSans 448 90 0 0 la_data_out[104]
port 276 nsew signal tristate
flabel metal2 s 499366 -960 499478 480 0 FreeSans 448 90 0 0 la_data_out[105]
port 277 nsew signal tristate
flabel metal2 s 502954 -960 503066 480 0 FreeSans 448 90 0 0 la_data_out[106]
port 278 nsew signal tristate
flabel metal2 s 506450 -960 506562 480 0 FreeSans 448 90 0 0 la_data_out[107]
port 279 nsew signal tristate
flabel metal2 s 510038 -960 510150 480 0 FreeSans 448 90 0 0 la_data_out[108]
port 280 nsew signal tristate
flabel metal2 s 513534 -960 513646 480 0 FreeSans 448 90 0 0 la_data_out[109]
port 281 nsew signal tristate
flabel metal2 s 162462 -960 162574 480 0 FreeSans 448 90 0 0 la_data_out[10]
port 282 nsew signal tristate
flabel metal2 s 517122 -960 517234 480 0 FreeSans 448 90 0 0 la_data_out[110]
port 283 nsew signal tristate
flabel metal2 s 520710 -960 520822 480 0 FreeSans 448 90 0 0 la_data_out[111]
port 284 nsew signal tristate
flabel metal2 s 524206 -960 524318 480 0 FreeSans 448 90 0 0 la_data_out[112]
port 285 nsew signal tristate
flabel metal2 s 527794 -960 527906 480 0 FreeSans 448 90 0 0 la_data_out[113]
port 286 nsew signal tristate
flabel metal2 s 531290 -960 531402 480 0 FreeSans 448 90 0 0 la_data_out[114]
port 287 nsew signal tristate
flabel metal2 s 534878 -960 534990 480 0 FreeSans 448 90 0 0 la_data_out[115]
port 288 nsew signal tristate
flabel metal2 s 538374 -960 538486 480 0 FreeSans 448 90 0 0 la_data_out[116]
port 289 nsew signal tristate
flabel metal2 s 541962 -960 542074 480 0 FreeSans 448 90 0 0 la_data_out[117]
port 290 nsew signal tristate
flabel metal2 s 545458 -960 545570 480 0 FreeSans 448 90 0 0 la_data_out[118]
port 291 nsew signal tristate
flabel metal2 s 549046 -960 549158 480 0 FreeSans 448 90 0 0 la_data_out[119]
port 292 nsew signal tristate
flabel metal2 s 166050 -960 166162 480 0 FreeSans 448 90 0 0 la_data_out[11]
port 293 nsew signal tristate
flabel metal2 s 552634 -960 552746 480 0 FreeSans 448 90 0 0 la_data_out[120]
port 294 nsew signal tristate
flabel metal2 s 556130 -960 556242 480 0 FreeSans 448 90 0 0 la_data_out[121]
port 295 nsew signal tristate
flabel metal2 s 559718 -960 559830 480 0 FreeSans 448 90 0 0 la_data_out[122]
port 296 nsew signal tristate
flabel metal2 s 563214 -960 563326 480 0 FreeSans 448 90 0 0 la_data_out[123]
port 297 nsew signal tristate
flabel metal2 s 566802 -960 566914 480 0 FreeSans 448 90 0 0 la_data_out[124]
port 298 nsew signal tristate
flabel metal2 s 570298 -960 570410 480 0 FreeSans 448 90 0 0 la_data_out[125]
port 299 nsew signal tristate
flabel metal2 s 573886 -960 573998 480 0 FreeSans 448 90 0 0 la_data_out[126]
port 300 nsew signal tristate
flabel metal2 s 577382 -960 577494 480 0 FreeSans 448 90 0 0 la_data_out[127]
port 301 nsew signal tristate
flabel metal2 s 169546 -960 169658 480 0 FreeSans 448 90 0 0 la_data_out[12]
port 302 nsew signal tristate
flabel metal2 s 173134 -960 173246 480 0 FreeSans 448 90 0 0 la_data_out[13]
port 303 nsew signal tristate
flabel metal2 s 176630 -960 176742 480 0 FreeSans 448 90 0 0 la_data_out[14]
port 304 nsew signal tristate
flabel metal2 s 180218 -960 180330 480 0 FreeSans 448 90 0 0 la_data_out[15]
port 305 nsew signal tristate
flabel metal2 s 183714 -960 183826 480 0 FreeSans 448 90 0 0 la_data_out[16]
port 306 nsew signal tristate
flabel metal2 s 187302 -960 187414 480 0 FreeSans 448 90 0 0 la_data_out[17]
port 307 nsew signal tristate
flabel metal2 s 190798 -960 190910 480 0 FreeSans 448 90 0 0 la_data_out[18]
port 308 nsew signal tristate
flabel metal2 s 194386 -960 194498 480 0 FreeSans 448 90 0 0 la_data_out[19]
port 309 nsew signal tristate
flabel metal2 s 130538 -960 130650 480 0 FreeSans 448 90 0 0 la_data_out[1]
port 310 nsew signal tristate
flabel metal2 s 197882 -960 197994 480 0 FreeSans 448 90 0 0 la_data_out[20]
port 311 nsew signal tristate
flabel metal2 s 201470 -960 201582 480 0 FreeSans 448 90 0 0 la_data_out[21]
port 312 nsew signal tristate
flabel metal2 s 205058 -960 205170 480 0 FreeSans 448 90 0 0 la_data_out[22]
port 313 nsew signal tristate
flabel metal2 s 208554 -960 208666 480 0 FreeSans 448 90 0 0 la_data_out[23]
port 314 nsew signal tristate
flabel metal2 s 212142 -960 212254 480 0 FreeSans 448 90 0 0 la_data_out[24]
port 315 nsew signal tristate
flabel metal2 s 215638 -960 215750 480 0 FreeSans 448 90 0 0 la_data_out[25]
port 316 nsew signal tristate
flabel metal2 s 219226 -960 219338 480 0 FreeSans 448 90 0 0 la_data_out[26]
port 317 nsew signal tristate
flabel metal2 s 222722 -960 222834 480 0 FreeSans 448 90 0 0 la_data_out[27]
port 318 nsew signal tristate
flabel metal2 s 226310 -960 226422 480 0 FreeSans 448 90 0 0 la_data_out[28]
port 319 nsew signal tristate
flabel metal2 s 229806 -960 229918 480 0 FreeSans 448 90 0 0 la_data_out[29]
port 320 nsew signal tristate
flabel metal2 s 134126 -960 134238 480 0 FreeSans 448 90 0 0 la_data_out[2]
port 321 nsew signal tristate
flabel metal2 s 233394 -960 233506 480 0 FreeSans 448 90 0 0 la_data_out[30]
port 322 nsew signal tristate
flabel metal2 s 236982 -960 237094 480 0 FreeSans 448 90 0 0 la_data_out[31]
port 323 nsew signal tristate
flabel metal2 s 240478 -960 240590 480 0 FreeSans 448 90 0 0 la_data_out[32]
port 324 nsew signal tristate
flabel metal2 s 244066 -960 244178 480 0 FreeSans 448 90 0 0 la_data_out[33]
port 325 nsew signal tristate
flabel metal2 s 247562 -960 247674 480 0 FreeSans 448 90 0 0 la_data_out[34]
port 326 nsew signal tristate
flabel metal2 s 251150 -960 251262 480 0 FreeSans 448 90 0 0 la_data_out[35]
port 327 nsew signal tristate
flabel metal2 s 254646 -960 254758 480 0 FreeSans 448 90 0 0 la_data_out[36]
port 328 nsew signal tristate
flabel metal2 s 258234 -960 258346 480 0 FreeSans 448 90 0 0 la_data_out[37]
port 329 nsew signal tristate
flabel metal2 s 261730 -960 261842 480 0 FreeSans 448 90 0 0 la_data_out[38]
port 330 nsew signal tristate
flabel metal2 s 265318 -960 265430 480 0 FreeSans 448 90 0 0 la_data_out[39]
port 331 nsew signal tristate
flabel metal2 s 137622 -960 137734 480 0 FreeSans 448 90 0 0 la_data_out[3]
port 332 nsew signal tristate
flabel metal2 s 268814 -960 268926 480 0 FreeSans 448 90 0 0 la_data_out[40]
port 333 nsew signal tristate
flabel metal2 s 272402 -960 272514 480 0 FreeSans 448 90 0 0 la_data_out[41]
port 334 nsew signal tristate
flabel metal2 s 275990 -960 276102 480 0 FreeSans 448 90 0 0 la_data_out[42]
port 335 nsew signal tristate
flabel metal2 s 279486 -960 279598 480 0 FreeSans 448 90 0 0 la_data_out[43]
port 336 nsew signal tristate
flabel metal2 s 283074 -960 283186 480 0 FreeSans 448 90 0 0 la_data_out[44]
port 337 nsew signal tristate
flabel metal2 s 286570 -960 286682 480 0 FreeSans 448 90 0 0 la_data_out[45]
port 338 nsew signal tristate
flabel metal2 s 290158 -960 290270 480 0 FreeSans 448 90 0 0 la_data_out[46]
port 339 nsew signal tristate
flabel metal2 s 293654 -960 293766 480 0 FreeSans 448 90 0 0 la_data_out[47]
port 340 nsew signal tristate
flabel metal2 s 297242 -960 297354 480 0 FreeSans 448 90 0 0 la_data_out[48]
port 341 nsew signal tristate
flabel metal2 s 300738 -960 300850 480 0 FreeSans 448 90 0 0 la_data_out[49]
port 342 nsew signal tristate
flabel metal2 s 141210 -960 141322 480 0 FreeSans 448 90 0 0 la_data_out[4]
port 343 nsew signal tristate
flabel metal2 s 304326 -960 304438 480 0 FreeSans 448 90 0 0 la_data_out[50]
port 344 nsew signal tristate
flabel metal2 s 307914 -960 308026 480 0 FreeSans 448 90 0 0 la_data_out[51]
port 345 nsew signal tristate
flabel metal2 s 311410 -960 311522 480 0 FreeSans 448 90 0 0 la_data_out[52]
port 346 nsew signal tristate
flabel metal2 s 314998 -960 315110 480 0 FreeSans 448 90 0 0 la_data_out[53]
port 347 nsew signal tristate
flabel metal2 s 318494 -960 318606 480 0 FreeSans 448 90 0 0 la_data_out[54]
port 348 nsew signal tristate
flabel metal2 s 322082 -960 322194 480 0 FreeSans 448 90 0 0 la_data_out[55]
port 349 nsew signal tristate
flabel metal2 s 325578 -960 325690 480 0 FreeSans 448 90 0 0 la_data_out[56]
port 350 nsew signal tristate
flabel metal2 s 329166 -960 329278 480 0 FreeSans 448 90 0 0 la_data_out[57]
port 351 nsew signal tristate
flabel metal2 s 332662 -960 332774 480 0 FreeSans 448 90 0 0 la_data_out[58]
port 352 nsew signal tristate
flabel metal2 s 336250 -960 336362 480 0 FreeSans 448 90 0 0 la_data_out[59]
port 353 nsew signal tristate
flabel metal2 s 144706 -960 144818 480 0 FreeSans 448 90 0 0 la_data_out[5]
port 354 nsew signal tristate
flabel metal2 s 339838 -960 339950 480 0 FreeSans 448 90 0 0 la_data_out[60]
port 355 nsew signal tristate
flabel metal2 s 343334 -960 343446 480 0 FreeSans 448 90 0 0 la_data_out[61]
port 356 nsew signal tristate
flabel metal2 s 346922 -960 347034 480 0 FreeSans 448 90 0 0 la_data_out[62]
port 357 nsew signal tristate
flabel metal2 s 350418 -960 350530 480 0 FreeSans 448 90 0 0 la_data_out[63]
port 358 nsew signal tristate
flabel metal2 s 354006 -960 354118 480 0 FreeSans 448 90 0 0 la_data_out[64]
port 359 nsew signal tristate
flabel metal2 s 357502 -960 357614 480 0 FreeSans 448 90 0 0 la_data_out[65]
port 360 nsew signal tristate
flabel metal2 s 361090 -960 361202 480 0 FreeSans 448 90 0 0 la_data_out[66]
port 361 nsew signal tristate
flabel metal2 s 364586 -960 364698 480 0 FreeSans 448 90 0 0 la_data_out[67]
port 362 nsew signal tristate
flabel metal2 s 368174 -960 368286 480 0 FreeSans 448 90 0 0 la_data_out[68]
port 363 nsew signal tristate
flabel metal2 s 371670 -960 371782 480 0 FreeSans 448 90 0 0 la_data_out[69]
port 364 nsew signal tristate
flabel metal2 s 148294 -960 148406 480 0 FreeSans 448 90 0 0 la_data_out[6]
port 365 nsew signal tristate
flabel metal2 s 375258 -960 375370 480 0 FreeSans 448 90 0 0 la_data_out[70]
port 366 nsew signal tristate
flabel metal2 s 378846 -960 378958 480 0 FreeSans 448 90 0 0 la_data_out[71]
port 367 nsew signal tristate
flabel metal2 s 382342 -960 382454 480 0 FreeSans 448 90 0 0 la_data_out[72]
port 368 nsew signal tristate
flabel metal2 s 385930 -960 386042 480 0 FreeSans 448 90 0 0 la_data_out[73]
port 369 nsew signal tristate
flabel metal2 s 389426 -960 389538 480 0 FreeSans 448 90 0 0 la_data_out[74]
port 370 nsew signal tristate
flabel metal2 s 393014 -960 393126 480 0 FreeSans 448 90 0 0 la_data_out[75]
port 371 nsew signal tristate
flabel metal2 s 396510 -960 396622 480 0 FreeSans 448 90 0 0 la_data_out[76]
port 372 nsew signal tristate
flabel metal2 s 400098 -960 400210 480 0 FreeSans 448 90 0 0 la_data_out[77]
port 373 nsew signal tristate
flabel metal2 s 403594 -960 403706 480 0 FreeSans 448 90 0 0 la_data_out[78]
port 374 nsew signal tristate
flabel metal2 s 407182 -960 407294 480 0 FreeSans 448 90 0 0 la_data_out[79]
port 375 nsew signal tristate
flabel metal2 s 151790 -960 151902 480 0 FreeSans 448 90 0 0 la_data_out[7]
port 376 nsew signal tristate
flabel metal2 s 410770 -960 410882 480 0 FreeSans 448 90 0 0 la_data_out[80]
port 377 nsew signal tristate
flabel metal2 s 414266 -960 414378 480 0 FreeSans 448 90 0 0 la_data_out[81]
port 378 nsew signal tristate
flabel metal2 s 417854 -960 417966 480 0 FreeSans 448 90 0 0 la_data_out[82]
port 379 nsew signal tristate
flabel metal2 s 421350 -960 421462 480 0 FreeSans 448 90 0 0 la_data_out[83]
port 380 nsew signal tristate
flabel metal2 s 424938 -960 425050 480 0 FreeSans 448 90 0 0 la_data_out[84]
port 381 nsew signal tristate
flabel metal2 s 428434 -960 428546 480 0 FreeSans 448 90 0 0 la_data_out[85]
port 382 nsew signal tristate
flabel metal2 s 432022 -960 432134 480 0 FreeSans 448 90 0 0 la_data_out[86]
port 383 nsew signal tristate
flabel metal2 s 435518 -960 435630 480 0 FreeSans 448 90 0 0 la_data_out[87]
port 384 nsew signal tristate
flabel metal2 s 439106 -960 439218 480 0 FreeSans 448 90 0 0 la_data_out[88]
port 385 nsew signal tristate
flabel metal2 s 442602 -960 442714 480 0 FreeSans 448 90 0 0 la_data_out[89]
port 386 nsew signal tristate
flabel metal2 s 155378 -960 155490 480 0 FreeSans 448 90 0 0 la_data_out[8]
port 387 nsew signal tristate
flabel metal2 s 446190 -960 446302 480 0 FreeSans 448 90 0 0 la_data_out[90]
port 388 nsew signal tristate
flabel metal2 s 449778 -960 449890 480 0 FreeSans 448 90 0 0 la_data_out[91]
port 389 nsew signal tristate
flabel metal2 s 453274 -960 453386 480 0 FreeSans 448 90 0 0 la_data_out[92]
port 390 nsew signal tristate
flabel metal2 s 456862 -960 456974 480 0 FreeSans 448 90 0 0 la_data_out[93]
port 391 nsew signal tristate
flabel metal2 s 460358 -960 460470 480 0 FreeSans 448 90 0 0 la_data_out[94]
port 392 nsew signal tristate
flabel metal2 s 463946 -960 464058 480 0 FreeSans 448 90 0 0 la_data_out[95]
port 393 nsew signal tristate
flabel metal2 s 467442 -960 467554 480 0 FreeSans 448 90 0 0 la_data_out[96]
port 394 nsew signal tristate
flabel metal2 s 471030 -960 471142 480 0 FreeSans 448 90 0 0 la_data_out[97]
port 395 nsew signal tristate
flabel metal2 s 474526 -960 474638 480 0 FreeSans 448 90 0 0 la_data_out[98]
port 396 nsew signal tristate
flabel metal2 s 478114 -960 478226 480 0 FreeSans 448 90 0 0 la_data_out[99]
port 397 nsew signal tristate
flabel metal2 s 158874 -960 158986 480 0 FreeSans 448 90 0 0 la_data_out[9]
port 398 nsew signal tristate
flabel metal2 s 128146 -960 128258 480 0 FreeSans 448 90 0 0 la_oenb[0]
port 399 nsew signal input
flabel metal2 s 482806 -960 482918 480 0 FreeSans 448 90 0 0 la_oenb[100]
port 400 nsew signal input
flabel metal2 s 486394 -960 486506 480 0 FreeSans 448 90 0 0 la_oenb[101]
port 401 nsew signal input
flabel metal2 s 489890 -960 490002 480 0 FreeSans 448 90 0 0 la_oenb[102]
port 402 nsew signal input
flabel metal2 s 493478 -960 493590 480 0 FreeSans 448 90 0 0 la_oenb[103]
port 403 nsew signal input
flabel metal2 s 497066 -960 497178 480 0 FreeSans 448 90 0 0 la_oenb[104]
port 404 nsew signal input
flabel metal2 s 500562 -960 500674 480 0 FreeSans 448 90 0 0 la_oenb[105]
port 405 nsew signal input
flabel metal2 s 504150 -960 504262 480 0 FreeSans 448 90 0 0 la_oenb[106]
port 406 nsew signal input
flabel metal2 s 507646 -960 507758 480 0 FreeSans 448 90 0 0 la_oenb[107]
port 407 nsew signal input
flabel metal2 s 511234 -960 511346 480 0 FreeSans 448 90 0 0 la_oenb[108]
port 408 nsew signal input
flabel metal2 s 514730 -960 514842 480 0 FreeSans 448 90 0 0 la_oenb[109]
port 409 nsew signal input
flabel metal2 s 163658 -960 163770 480 0 FreeSans 448 90 0 0 la_oenb[10]
port 410 nsew signal input
flabel metal2 s 518318 -960 518430 480 0 FreeSans 448 90 0 0 la_oenb[110]
port 411 nsew signal input
flabel metal2 s 521814 -960 521926 480 0 FreeSans 448 90 0 0 la_oenb[111]
port 412 nsew signal input
flabel metal2 s 525402 -960 525514 480 0 FreeSans 448 90 0 0 la_oenb[112]
port 413 nsew signal input
flabel metal2 s 528990 -960 529102 480 0 FreeSans 448 90 0 0 la_oenb[113]
port 414 nsew signal input
flabel metal2 s 532486 -960 532598 480 0 FreeSans 448 90 0 0 la_oenb[114]
port 415 nsew signal input
flabel metal2 s 536074 -960 536186 480 0 FreeSans 448 90 0 0 la_oenb[115]
port 416 nsew signal input
flabel metal2 s 539570 -960 539682 480 0 FreeSans 448 90 0 0 la_oenb[116]
port 417 nsew signal input
flabel metal2 s 543158 -960 543270 480 0 FreeSans 448 90 0 0 la_oenb[117]
port 418 nsew signal input
flabel metal2 s 546654 -960 546766 480 0 FreeSans 448 90 0 0 la_oenb[118]
port 419 nsew signal input
flabel metal2 s 550242 -960 550354 480 0 FreeSans 448 90 0 0 la_oenb[119]
port 420 nsew signal input
flabel metal2 s 167154 -960 167266 480 0 FreeSans 448 90 0 0 la_oenb[11]
port 421 nsew signal input
flabel metal2 s 553738 -960 553850 480 0 FreeSans 448 90 0 0 la_oenb[120]
port 422 nsew signal input
flabel metal2 s 557326 -960 557438 480 0 FreeSans 448 90 0 0 la_oenb[121]
port 423 nsew signal input
flabel metal2 s 560822 -960 560934 480 0 FreeSans 448 90 0 0 la_oenb[122]
port 424 nsew signal input
flabel metal2 s 564410 -960 564522 480 0 FreeSans 448 90 0 0 la_oenb[123]
port 425 nsew signal input
flabel metal2 s 567998 -960 568110 480 0 FreeSans 448 90 0 0 la_oenb[124]
port 426 nsew signal input
flabel metal2 s 571494 -960 571606 480 0 FreeSans 448 90 0 0 la_oenb[125]
port 427 nsew signal input
flabel metal2 s 575082 -960 575194 480 0 FreeSans 448 90 0 0 la_oenb[126]
port 428 nsew signal input
flabel metal2 s 578578 -960 578690 480 0 FreeSans 448 90 0 0 la_oenb[127]
port 429 nsew signal input
flabel metal2 s 170742 -960 170854 480 0 FreeSans 448 90 0 0 la_oenb[12]
port 430 nsew signal input
flabel metal2 s 174238 -960 174350 480 0 FreeSans 448 90 0 0 la_oenb[13]
port 431 nsew signal input
flabel metal2 s 177826 -960 177938 480 0 FreeSans 448 90 0 0 la_oenb[14]
port 432 nsew signal input
flabel metal2 s 181414 -960 181526 480 0 FreeSans 448 90 0 0 la_oenb[15]
port 433 nsew signal input
flabel metal2 s 184910 -960 185022 480 0 FreeSans 448 90 0 0 la_oenb[16]
port 434 nsew signal input
flabel metal2 s 188498 -960 188610 480 0 FreeSans 448 90 0 0 la_oenb[17]
port 435 nsew signal input
flabel metal2 s 191994 -960 192106 480 0 FreeSans 448 90 0 0 la_oenb[18]
port 436 nsew signal input
flabel metal2 s 195582 -960 195694 480 0 FreeSans 448 90 0 0 la_oenb[19]
port 437 nsew signal input
flabel metal2 s 131734 -960 131846 480 0 FreeSans 448 90 0 0 la_oenb[1]
port 438 nsew signal input
flabel metal2 s 199078 -960 199190 480 0 FreeSans 448 90 0 0 la_oenb[20]
port 439 nsew signal input
flabel metal2 s 202666 -960 202778 480 0 FreeSans 448 90 0 0 la_oenb[21]
port 440 nsew signal input
flabel metal2 s 206162 -960 206274 480 0 FreeSans 448 90 0 0 la_oenb[22]
port 441 nsew signal input
flabel metal2 s 209750 -960 209862 480 0 FreeSans 448 90 0 0 la_oenb[23]
port 442 nsew signal input
flabel metal2 s 213338 -960 213450 480 0 FreeSans 448 90 0 0 la_oenb[24]
port 443 nsew signal input
flabel metal2 s 216834 -960 216946 480 0 FreeSans 448 90 0 0 la_oenb[25]
port 444 nsew signal input
flabel metal2 s 220422 -960 220534 480 0 FreeSans 448 90 0 0 la_oenb[26]
port 445 nsew signal input
flabel metal2 s 223918 -960 224030 480 0 FreeSans 448 90 0 0 la_oenb[27]
port 446 nsew signal input
flabel metal2 s 227506 -960 227618 480 0 FreeSans 448 90 0 0 la_oenb[28]
port 447 nsew signal input
flabel metal2 s 231002 -960 231114 480 0 FreeSans 448 90 0 0 la_oenb[29]
port 448 nsew signal input
flabel metal2 s 135230 -960 135342 480 0 FreeSans 448 90 0 0 la_oenb[2]
port 449 nsew signal input
flabel metal2 s 234590 -960 234702 480 0 FreeSans 448 90 0 0 la_oenb[30]
port 450 nsew signal input
flabel metal2 s 238086 -960 238198 480 0 FreeSans 448 90 0 0 la_oenb[31]
port 451 nsew signal input
flabel metal2 s 241674 -960 241786 480 0 FreeSans 448 90 0 0 la_oenb[32]
port 452 nsew signal input
flabel metal2 s 245170 -960 245282 480 0 FreeSans 448 90 0 0 la_oenb[33]
port 453 nsew signal input
flabel metal2 s 248758 -960 248870 480 0 FreeSans 448 90 0 0 la_oenb[34]
port 454 nsew signal input
flabel metal2 s 252346 -960 252458 480 0 FreeSans 448 90 0 0 la_oenb[35]
port 455 nsew signal input
flabel metal2 s 255842 -960 255954 480 0 FreeSans 448 90 0 0 la_oenb[36]
port 456 nsew signal input
flabel metal2 s 259430 -960 259542 480 0 FreeSans 448 90 0 0 la_oenb[37]
port 457 nsew signal input
flabel metal2 s 262926 -960 263038 480 0 FreeSans 448 90 0 0 la_oenb[38]
port 458 nsew signal input
flabel metal2 s 266514 -960 266626 480 0 FreeSans 448 90 0 0 la_oenb[39]
port 459 nsew signal input
flabel metal2 s 138818 -960 138930 480 0 FreeSans 448 90 0 0 la_oenb[3]
port 460 nsew signal input
flabel metal2 s 270010 -960 270122 480 0 FreeSans 448 90 0 0 la_oenb[40]
port 461 nsew signal input
flabel metal2 s 273598 -960 273710 480 0 FreeSans 448 90 0 0 la_oenb[41]
port 462 nsew signal input
flabel metal2 s 277094 -960 277206 480 0 FreeSans 448 90 0 0 la_oenb[42]
port 463 nsew signal input
flabel metal2 s 280682 -960 280794 480 0 FreeSans 448 90 0 0 la_oenb[43]
port 464 nsew signal input
flabel metal2 s 284270 -960 284382 480 0 FreeSans 448 90 0 0 la_oenb[44]
port 465 nsew signal input
flabel metal2 s 287766 -960 287878 480 0 FreeSans 448 90 0 0 la_oenb[45]
port 466 nsew signal input
flabel metal2 s 291354 -960 291466 480 0 FreeSans 448 90 0 0 la_oenb[46]
port 467 nsew signal input
flabel metal2 s 294850 -960 294962 480 0 FreeSans 448 90 0 0 la_oenb[47]
port 468 nsew signal input
flabel metal2 s 298438 -960 298550 480 0 FreeSans 448 90 0 0 la_oenb[48]
port 469 nsew signal input
flabel metal2 s 301934 -960 302046 480 0 FreeSans 448 90 0 0 la_oenb[49]
port 470 nsew signal input
flabel metal2 s 142406 -960 142518 480 0 FreeSans 448 90 0 0 la_oenb[4]
port 471 nsew signal input
flabel metal2 s 305522 -960 305634 480 0 FreeSans 448 90 0 0 la_oenb[50]
port 472 nsew signal input
flabel metal2 s 309018 -960 309130 480 0 FreeSans 448 90 0 0 la_oenb[51]
port 473 nsew signal input
flabel metal2 s 312606 -960 312718 480 0 FreeSans 448 90 0 0 la_oenb[52]
port 474 nsew signal input
flabel metal2 s 316194 -960 316306 480 0 FreeSans 448 90 0 0 la_oenb[53]
port 475 nsew signal input
flabel metal2 s 319690 -960 319802 480 0 FreeSans 448 90 0 0 la_oenb[54]
port 476 nsew signal input
flabel metal2 s 323278 -960 323390 480 0 FreeSans 448 90 0 0 la_oenb[55]
port 477 nsew signal input
flabel metal2 s 326774 -960 326886 480 0 FreeSans 448 90 0 0 la_oenb[56]
port 478 nsew signal input
flabel metal2 s 330362 -960 330474 480 0 FreeSans 448 90 0 0 la_oenb[57]
port 479 nsew signal input
flabel metal2 s 333858 -960 333970 480 0 FreeSans 448 90 0 0 la_oenb[58]
port 480 nsew signal input
flabel metal2 s 337446 -960 337558 480 0 FreeSans 448 90 0 0 la_oenb[59]
port 481 nsew signal input
flabel metal2 s 145902 -960 146014 480 0 FreeSans 448 90 0 0 la_oenb[5]
port 482 nsew signal input
flabel metal2 s 340942 -960 341054 480 0 FreeSans 448 90 0 0 la_oenb[60]
port 483 nsew signal input
flabel metal2 s 344530 -960 344642 480 0 FreeSans 448 90 0 0 la_oenb[61]
port 484 nsew signal input
flabel metal2 s 348026 -960 348138 480 0 FreeSans 448 90 0 0 la_oenb[62]
port 485 nsew signal input
flabel metal2 s 351614 -960 351726 480 0 FreeSans 448 90 0 0 la_oenb[63]
port 486 nsew signal input
flabel metal2 s 355202 -960 355314 480 0 FreeSans 448 90 0 0 la_oenb[64]
port 487 nsew signal input
flabel metal2 s 358698 -960 358810 480 0 FreeSans 448 90 0 0 la_oenb[65]
port 488 nsew signal input
flabel metal2 s 362286 -960 362398 480 0 FreeSans 448 90 0 0 la_oenb[66]
port 489 nsew signal input
flabel metal2 s 365782 -960 365894 480 0 FreeSans 448 90 0 0 la_oenb[67]
port 490 nsew signal input
flabel metal2 s 369370 -960 369482 480 0 FreeSans 448 90 0 0 la_oenb[68]
port 491 nsew signal input
flabel metal2 s 372866 -960 372978 480 0 FreeSans 448 90 0 0 la_oenb[69]
port 492 nsew signal input
flabel metal2 s 149490 -960 149602 480 0 FreeSans 448 90 0 0 la_oenb[6]
port 493 nsew signal input
flabel metal2 s 376454 -960 376566 480 0 FreeSans 448 90 0 0 la_oenb[70]
port 494 nsew signal input
flabel metal2 s 379950 -960 380062 480 0 FreeSans 448 90 0 0 la_oenb[71]
port 495 nsew signal input
flabel metal2 s 383538 -960 383650 480 0 FreeSans 448 90 0 0 la_oenb[72]
port 496 nsew signal input
flabel metal2 s 387126 -960 387238 480 0 FreeSans 448 90 0 0 la_oenb[73]
port 497 nsew signal input
flabel metal2 s 390622 -960 390734 480 0 FreeSans 448 90 0 0 la_oenb[74]
port 498 nsew signal input
flabel metal2 s 394210 -960 394322 480 0 FreeSans 448 90 0 0 la_oenb[75]
port 499 nsew signal input
flabel metal2 s 397706 -960 397818 480 0 FreeSans 448 90 0 0 la_oenb[76]
port 500 nsew signal input
flabel metal2 s 401294 -960 401406 480 0 FreeSans 448 90 0 0 la_oenb[77]
port 501 nsew signal input
flabel metal2 s 404790 -960 404902 480 0 FreeSans 448 90 0 0 la_oenb[78]
port 502 nsew signal input
flabel metal2 s 408378 -960 408490 480 0 FreeSans 448 90 0 0 la_oenb[79]
port 503 nsew signal input
flabel metal2 s 152986 -960 153098 480 0 FreeSans 448 90 0 0 la_oenb[7]
port 504 nsew signal input
flabel metal2 s 411874 -960 411986 480 0 FreeSans 448 90 0 0 la_oenb[80]
port 505 nsew signal input
flabel metal2 s 415462 -960 415574 480 0 FreeSans 448 90 0 0 la_oenb[81]
port 506 nsew signal input
flabel metal2 s 418958 -960 419070 480 0 FreeSans 448 90 0 0 la_oenb[82]
port 507 nsew signal input
flabel metal2 s 422546 -960 422658 480 0 FreeSans 448 90 0 0 la_oenb[83]
port 508 nsew signal input
flabel metal2 s 426134 -960 426246 480 0 FreeSans 448 90 0 0 la_oenb[84]
port 509 nsew signal input
flabel metal2 s 429630 -960 429742 480 0 FreeSans 448 90 0 0 la_oenb[85]
port 510 nsew signal input
flabel metal2 s 433218 -960 433330 480 0 FreeSans 448 90 0 0 la_oenb[86]
port 511 nsew signal input
flabel metal2 s 436714 -960 436826 480 0 FreeSans 448 90 0 0 la_oenb[87]
port 512 nsew signal input
flabel metal2 s 440302 -960 440414 480 0 FreeSans 448 90 0 0 la_oenb[88]
port 513 nsew signal input
flabel metal2 s 443798 -960 443910 480 0 FreeSans 448 90 0 0 la_oenb[89]
port 514 nsew signal input
flabel metal2 s 156574 -960 156686 480 0 FreeSans 448 90 0 0 la_oenb[8]
port 515 nsew signal input
flabel metal2 s 447386 -960 447498 480 0 FreeSans 448 90 0 0 la_oenb[90]
port 516 nsew signal input
flabel metal2 s 450882 -960 450994 480 0 FreeSans 448 90 0 0 la_oenb[91]
port 517 nsew signal input
flabel metal2 s 454470 -960 454582 480 0 FreeSans 448 90 0 0 la_oenb[92]
port 518 nsew signal input
flabel metal2 s 458058 -960 458170 480 0 FreeSans 448 90 0 0 la_oenb[93]
port 519 nsew signal input
flabel metal2 s 461554 -960 461666 480 0 FreeSans 448 90 0 0 la_oenb[94]
port 520 nsew signal input
flabel metal2 s 465142 -960 465254 480 0 FreeSans 448 90 0 0 la_oenb[95]
port 521 nsew signal input
flabel metal2 s 468638 -960 468750 480 0 FreeSans 448 90 0 0 la_oenb[96]
port 522 nsew signal input
flabel metal2 s 472226 -960 472338 480 0 FreeSans 448 90 0 0 la_oenb[97]
port 523 nsew signal input
flabel metal2 s 475722 -960 475834 480 0 FreeSans 448 90 0 0 la_oenb[98]
port 524 nsew signal input
flabel metal2 s 479310 -960 479422 480 0 FreeSans 448 90 0 0 la_oenb[99]
port 525 nsew signal input
flabel metal2 s 160070 -960 160182 480 0 FreeSans 448 90 0 0 la_oenb[9]
port 526 nsew signal input
flabel metal2 s 579774 -960 579886 480 0 FreeSans 448 90 0 0 user_clock2
port 527 nsew signal input
flabel metal2 s 580970 -960 581082 480 0 FreeSans 448 90 0 0 user_irq[0]
port 528 nsew signal tristate
flabel metal2 s 582166 -960 582278 480 0 FreeSans 448 90 0 0 user_irq[1]
port 529 nsew signal tristate
flabel metal2 s 583362 -960 583474 480 0 FreeSans 448 90 0 0 user_irq[2]
port 530 nsew signal tristate
flabel metal4 s -2006 -934 -1386 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 -934 585930 -314 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 704250 585930 704870 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 585310 -934 585930 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 1794 -7654 2414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 37794 -7654 38414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 73794 -7654 74414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 109794 -7654 110414 498000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 109794 591292 110414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 145794 -7654 146414 498000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 145794 591292 146414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 181794 -7654 182414 498000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 181794 591292 182414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 217794 -7654 218414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 253794 -7654 254414 336000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 253794 384000 254414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 289794 -7654 290414 98000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 289794 158000 290414 336000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 289794 384000 290414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 325794 -7654 326414 98000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 325794 158000 326414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 361794 -7654 362414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 397794 -7654 398414 498000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 397794 591292 398414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 433794 -7654 434414 498000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 433794 591292 434414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 469794 -7654 470414 498000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 469794 591292 470414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 505794 -7654 506414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 541794 -7654 542414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 577794 -7654 578414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 2866 592650 3486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 38866 592650 39486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 74866 592650 75486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 110866 592650 111486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 146866 592650 147486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 182866 592650 183486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 218866 592650 219486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 254866 592650 255486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 290866 592650 291486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 326866 592650 327486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 362866 592650 363486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 398866 592650 399486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 434866 592650 435486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 470866 592650 471486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 506866 592650 507486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 542866 592650 543486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 578866 592650 579486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 614866 592650 615486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 650866 592650 651486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 686866 592650 687486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s -3926 -2854 -3306 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 -2854 587850 -2234 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 706170 587850 706790 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 587230 -2854 587850 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 10794 -7654 11414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 46794 -7654 47414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 82794 -7654 83414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 118794 -7654 119414 498000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 118794 591292 119414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 154794 -7654 155414 498000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 154794 591292 155414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 190794 -7654 191414 498000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 190794 591292 191414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 226794 -7654 227414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 262794 -7654 263414 98000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 262794 158000 263414 336000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 262794 384000 263414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 298794 -7654 299414 98000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 298794 158000 299414 336000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 298794 384000 299414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 334794 -7654 335414 98000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 334794 158000 335414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 370794 -7654 371414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 406794 -7654 407414 498000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 406794 591292 407414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 442794 -7654 443414 498000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 442794 591292 443414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 478794 -7654 479414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 514794 -7654 515414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 550794 -7654 551414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 11866 592650 12486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 47866 592650 48486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 83866 592650 84486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 119866 592650 120486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 155866 592650 156486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 191866 592650 192486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 227866 592650 228486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 263866 592650 264486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 299866 592650 300486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 335866 592650 336486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 371866 592650 372486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 407866 592650 408486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 443866 592650 444486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 479866 592650 480486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 515866 592650 516486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 551866 592650 552486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 587866 592650 588486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 623866 592650 624486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 659866 592650 660486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 695866 592650 696486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s -5846 -4774 -5226 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 -4774 589770 -4154 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 708090 589770 708710 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 589150 -4774 589770 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 19794 -7654 20414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 55794 -7654 56414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 91794 -7654 92414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 127794 -7654 128414 498000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 127794 591292 128414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 163794 -7654 164414 498000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 163794 591292 164414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 199794 -7654 200414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 235794 -7654 236414 336000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 235794 384000 236414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 271794 -7654 272414 98000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 271794 158000 272414 336000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 271794 384000 272414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 307794 -7654 308414 98000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 307794 158000 308414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 343794 -7654 344414 98000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 343794 158000 344414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 379794 -7654 380414 498000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 379794 591292 380414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 415794 -7654 416414 498000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 415794 591292 416414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 451794 -7654 452414 498000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 451794 591292 452414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 487794 -7654 488414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 523794 -7654 524414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 559794 -7654 560414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 20866 592650 21486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 56866 592650 57486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 92866 592650 93486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 128866 592650 129486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 164866 592650 165486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 200866 592650 201486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 236866 592650 237486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 272866 592650 273486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 308866 592650 309486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 344866 592650 345486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 380866 592650 381486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 416866 592650 417486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 452866 592650 453486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 488866 592650 489486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 524866 592650 525486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 560866 592650 561486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 596866 592650 597486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 632866 592650 633486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 668866 592650 669486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s -7766 -6694 -7146 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -7766 -6694 591690 -6074 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -7766 710010 591690 710630 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 591070 -6694 591690 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 28794 -7654 29414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 64794 -7654 65414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 100794 -7654 101414 498000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 100794 591292 101414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 136794 -7654 137414 498000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 136794 591292 137414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 172794 -7654 173414 498000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 172794 591292 173414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 208794 -7654 209414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 244794 -7654 245414 336000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 244794 384000 245414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 280794 -7654 281414 98000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 280794 158000 281414 336000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 280794 384000 281414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 316794 -7654 317414 98000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 316794 158000 317414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 352794 -7654 353414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 388794 -7654 389414 498000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 388794 591292 389414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 424794 -7654 425414 498000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 424794 591292 425414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 460794 -7654 461414 498000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 460794 591292 461414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 496794 -7654 497414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 532794 -7654 533414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 568794 -7654 569414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 29866 592650 30486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 65866 592650 66486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 101866 592650 102486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 137866 592650 138486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 173866 592650 174486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 209866 592650 210486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 245866 592650 246486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 281866 592650 282486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 317866 592650 318486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 353866 592650 354486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 389866 592650 390486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 425866 592650 426486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 461866 592650 462486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 497866 592650 498486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 533866 592650 534486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 569866 592650 570486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 605866 592650 606486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 641866 592650 642486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 677866 592650 678486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s -6806 -5734 -6186 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 -5734 590730 -5114 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 709050 590730 709670 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 590110 -5734 590730 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 24294 -7654 24914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 60294 -7654 60914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 96294 -7654 96914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 132294 -7654 132914 498000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 132294 591292 132914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 168294 -7654 168914 498000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 168294 591292 168914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 204294 -7654 204914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 240294 -7654 240914 336000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 240294 384000 240914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 276294 -7654 276914 98000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 276294 158000 276914 336000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 276294 384000 276914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 312294 -7654 312914 98000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 312294 158000 312914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 348294 -7654 348914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 384294 -7654 384914 498000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 384294 591292 384914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 420294 -7654 420914 498000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 420294 591292 420914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 456294 -7654 456914 498000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 456294 591292 456914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 492294 -7654 492914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 528294 -7654 528914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 564294 -7654 564914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 25366 592650 25986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 61366 592650 61986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 97366 592650 97986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 133366 592650 133986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 169366 592650 169986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 205366 592650 205986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 241366 592650 241986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 277366 592650 277986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 313366 592650 313986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 349366 592650 349986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 385366 592650 385986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 421366 592650 421986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 457366 592650 457986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 493366 592650 493986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 529366 592650 529986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 565366 592650 565986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 601366 592650 601986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 637366 592650 637986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 673366 592650 673986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s -8726 -7654 -8106 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 -7654 592650 -7034 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 710970 592650 711590 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 592030 -7654 592650 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 33294 -7654 33914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 69294 -7654 69914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 105294 -7654 105914 498000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 105294 591292 105914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 141294 -7654 141914 498000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 141294 591292 141914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 177294 -7654 177914 498000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 177294 591292 177914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 213294 -7654 213914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 249294 -7654 249914 336000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 249294 384000 249914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 285294 -7654 285914 98000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 285294 158000 285914 336000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 285294 384000 285914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 321294 -7654 321914 98000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 321294 158000 321914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 357294 -7654 357914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 393294 -7654 393914 498000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 393294 591292 393914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 429294 -7654 429914 498000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 429294 591292 429914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 465294 -7654 465914 498000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 465294 591292 465914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 501294 -7654 501914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 537294 -7654 537914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 573294 -7654 573914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 34366 592650 34986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 70366 592650 70986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 106366 592650 106986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 142366 592650 142986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 178366 592650 178986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 214366 592650 214986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 250366 592650 250986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 286366 592650 286986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 322366 592650 322986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 358366 592650 358986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 394366 592650 394986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 430366 592650 430986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 466366 592650 466986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 502366 592650 502986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 538366 592650 538986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 574366 592650 574986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 610366 592650 610986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 646366 592650 646986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 682366 592650 682986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s -2966 -1894 -2346 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 -1894 586890 -1274 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 705210 586890 705830 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 586270 -1894 586890 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 6294 -7654 6914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 42294 -7654 42914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 78294 -7654 78914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 114294 -7654 114914 498000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 114294 591292 114914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 150294 -7654 150914 498000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 150294 591292 150914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 186294 -7654 186914 498000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 186294 591292 186914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 222294 -7654 222914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 258294 -7654 258914 98000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 258294 158000 258914 336000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 258294 384000 258914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 294294 -7654 294914 98000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 294294 158000 294914 336000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 294294 384000 294914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 330294 -7654 330914 98000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 330294 158000 330914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 366294 -7654 366914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 402294 -7654 402914 498000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 402294 591292 402914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 438294 -7654 438914 498000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 438294 591292 438914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 474294 -7654 474914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 510294 -7654 510914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 546294 -7654 546914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 582294 -7654 582914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 7366 592650 7986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 43366 592650 43986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 79366 592650 79986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 115366 592650 115986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 151366 592650 151986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 187366 592650 187986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 223366 592650 223986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 259366 592650 259986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 295366 592650 295986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 331366 592650 331986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 367366 592650 367986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 403366 592650 403986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 439366 592650 439986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 475366 592650 475986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 511366 592650 511986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 547366 592650 547986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 583366 592650 583986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 619366 592650 619986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 655366 592650 655986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 691366 592650 691986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s -4886 -3814 -4266 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 -3814 588810 -3194 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 707130 588810 707750 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 588190 -3814 588810 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 15294 -7654 15914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 51294 -7654 51914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 87294 -7654 87914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 123294 -7654 123914 498000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 123294 591292 123914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 159294 -7654 159914 498000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 159294 591292 159914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 195294 -7654 195914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 231294 -7654 231914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 267294 -7654 267914 98000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 267294 158000 267914 336000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 267294 384000 267914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 303294 -7654 303914 98000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 303294 158000 303914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 339294 -7654 339914 98000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 339294 158000 339914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 375294 -7654 375914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 411294 -7654 411914 498000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 411294 591292 411914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 447294 -7654 447914 498000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 447294 591292 447914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 483294 -7654 483914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 519294 -7654 519914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 555294 -7654 555914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 16366 592650 16986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 52366 592650 52986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 88366 592650 88986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 124366 592650 124986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 160366 592650 160986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 196366 592650 196986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 232366 592650 232986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 268366 592650 268986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 304366 592650 304986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 340366 592650 340986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 376366 592650 376986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 412366 592650 412986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 448366 592650 448986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 484366 592650 484986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 520366 592650 520986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 556366 592650 556986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 592366 592650 592986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 628366 592650 628986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 664366 592650 664986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 700366 592650 700986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal2 s 542 -960 654 480 0 FreeSans 448 90 0 0 wb_clk_i
port 539 nsew signal input
flabel metal2 s 1646 -960 1758 480 0 FreeSans 448 90 0 0 wb_rst_i
port 540 nsew signal input
flabel metal2 s 2842 -960 2954 480 0 FreeSans 448 90 0 0 wbs_ack_o
port 541 nsew signal tristate
flabel metal2 s 7626 -960 7738 480 0 FreeSans 448 90 0 0 wbs_adr_i[0]
port 542 nsew signal input
flabel metal2 s 47830 -960 47942 480 0 FreeSans 448 90 0 0 wbs_adr_i[10]
port 543 nsew signal input
flabel metal2 s 51326 -960 51438 480 0 FreeSans 448 90 0 0 wbs_adr_i[11]
port 544 nsew signal input
flabel metal2 s 54914 -960 55026 480 0 FreeSans 448 90 0 0 wbs_adr_i[12]
port 545 nsew signal input
flabel metal2 s 58410 -960 58522 480 0 FreeSans 448 90 0 0 wbs_adr_i[13]
port 546 nsew signal input
flabel metal2 s 61998 -960 62110 480 0 FreeSans 448 90 0 0 wbs_adr_i[14]
port 547 nsew signal input
flabel metal2 s 65494 -960 65606 480 0 FreeSans 448 90 0 0 wbs_adr_i[15]
port 548 nsew signal input
flabel metal2 s 69082 -960 69194 480 0 FreeSans 448 90 0 0 wbs_adr_i[16]
port 549 nsew signal input
flabel metal2 s 72578 -960 72690 480 0 FreeSans 448 90 0 0 wbs_adr_i[17]
port 550 nsew signal input
flabel metal2 s 76166 -960 76278 480 0 FreeSans 448 90 0 0 wbs_adr_i[18]
port 551 nsew signal input
flabel metal2 s 79662 -960 79774 480 0 FreeSans 448 90 0 0 wbs_adr_i[19]
port 552 nsew signal input
flabel metal2 s 12318 -960 12430 480 0 FreeSans 448 90 0 0 wbs_adr_i[1]
port 553 nsew signal input
flabel metal2 s 83250 -960 83362 480 0 FreeSans 448 90 0 0 wbs_adr_i[20]
port 554 nsew signal input
flabel metal2 s 86838 -960 86950 480 0 FreeSans 448 90 0 0 wbs_adr_i[21]
port 555 nsew signal input
flabel metal2 s 90334 -960 90446 480 0 FreeSans 448 90 0 0 wbs_adr_i[22]
port 556 nsew signal input
flabel metal2 s 93922 -960 94034 480 0 FreeSans 448 90 0 0 wbs_adr_i[23]
port 557 nsew signal input
flabel metal2 s 97418 -960 97530 480 0 FreeSans 448 90 0 0 wbs_adr_i[24]
port 558 nsew signal input
flabel metal2 s 101006 -960 101118 480 0 FreeSans 448 90 0 0 wbs_adr_i[25]
port 559 nsew signal input
flabel metal2 s 104502 -960 104614 480 0 FreeSans 448 90 0 0 wbs_adr_i[26]
port 560 nsew signal input
flabel metal2 s 108090 -960 108202 480 0 FreeSans 448 90 0 0 wbs_adr_i[27]
port 561 nsew signal input
flabel metal2 s 111586 -960 111698 480 0 FreeSans 448 90 0 0 wbs_adr_i[28]
port 562 nsew signal input
flabel metal2 s 115174 -960 115286 480 0 FreeSans 448 90 0 0 wbs_adr_i[29]
port 563 nsew signal input
flabel metal2 s 17010 -960 17122 480 0 FreeSans 448 90 0 0 wbs_adr_i[2]
port 564 nsew signal input
flabel metal2 s 118762 -960 118874 480 0 FreeSans 448 90 0 0 wbs_adr_i[30]
port 565 nsew signal input
flabel metal2 s 122258 -960 122370 480 0 FreeSans 448 90 0 0 wbs_adr_i[31]
port 566 nsew signal input
flabel metal2 s 21794 -960 21906 480 0 FreeSans 448 90 0 0 wbs_adr_i[3]
port 567 nsew signal input
flabel metal2 s 26486 -960 26598 480 0 FreeSans 448 90 0 0 wbs_adr_i[4]
port 568 nsew signal input
flabel metal2 s 30074 -960 30186 480 0 FreeSans 448 90 0 0 wbs_adr_i[5]
port 569 nsew signal input
flabel metal2 s 33570 -960 33682 480 0 FreeSans 448 90 0 0 wbs_adr_i[6]
port 570 nsew signal input
flabel metal2 s 37158 -960 37270 480 0 FreeSans 448 90 0 0 wbs_adr_i[7]
port 571 nsew signal input
flabel metal2 s 40654 -960 40766 480 0 FreeSans 448 90 0 0 wbs_adr_i[8]
port 572 nsew signal input
flabel metal2 s 44242 -960 44354 480 0 FreeSans 448 90 0 0 wbs_adr_i[9]
port 573 nsew signal input
flabel metal2 s 4038 -960 4150 480 0 FreeSans 448 90 0 0 wbs_cyc_i
port 574 nsew signal input
flabel metal2 s 8730 -960 8842 480 0 FreeSans 448 90 0 0 wbs_dat_i[0]
port 575 nsew signal input
flabel metal2 s 48934 -960 49046 480 0 FreeSans 448 90 0 0 wbs_dat_i[10]
port 576 nsew signal input
flabel metal2 s 52522 -960 52634 480 0 FreeSans 448 90 0 0 wbs_dat_i[11]
port 577 nsew signal input
flabel metal2 s 56018 -960 56130 480 0 FreeSans 448 90 0 0 wbs_dat_i[12]
port 578 nsew signal input
flabel metal2 s 59606 -960 59718 480 0 FreeSans 448 90 0 0 wbs_dat_i[13]
port 579 nsew signal input
flabel metal2 s 63194 -960 63306 480 0 FreeSans 448 90 0 0 wbs_dat_i[14]
port 580 nsew signal input
flabel metal2 s 66690 -960 66802 480 0 FreeSans 448 90 0 0 wbs_dat_i[15]
port 581 nsew signal input
flabel metal2 s 70278 -960 70390 480 0 FreeSans 448 90 0 0 wbs_dat_i[16]
port 582 nsew signal input
flabel metal2 s 73774 -960 73886 480 0 FreeSans 448 90 0 0 wbs_dat_i[17]
port 583 nsew signal input
flabel metal2 s 77362 -960 77474 480 0 FreeSans 448 90 0 0 wbs_dat_i[18]
port 584 nsew signal input
flabel metal2 s 80858 -960 80970 480 0 FreeSans 448 90 0 0 wbs_dat_i[19]
port 585 nsew signal input
flabel metal2 s 13514 -960 13626 480 0 FreeSans 448 90 0 0 wbs_dat_i[1]
port 586 nsew signal input
flabel metal2 s 84446 -960 84558 480 0 FreeSans 448 90 0 0 wbs_dat_i[20]
port 587 nsew signal input
flabel metal2 s 87942 -960 88054 480 0 FreeSans 448 90 0 0 wbs_dat_i[21]
port 588 nsew signal input
flabel metal2 s 91530 -960 91642 480 0 FreeSans 448 90 0 0 wbs_dat_i[22]
port 589 nsew signal input
flabel metal2 s 95118 -960 95230 480 0 FreeSans 448 90 0 0 wbs_dat_i[23]
port 590 nsew signal input
flabel metal2 s 98614 -960 98726 480 0 FreeSans 448 90 0 0 wbs_dat_i[24]
port 591 nsew signal input
flabel metal2 s 102202 -960 102314 480 0 FreeSans 448 90 0 0 wbs_dat_i[25]
port 592 nsew signal input
flabel metal2 s 105698 -960 105810 480 0 FreeSans 448 90 0 0 wbs_dat_i[26]
port 593 nsew signal input
flabel metal2 s 109286 -960 109398 480 0 FreeSans 448 90 0 0 wbs_dat_i[27]
port 594 nsew signal input
flabel metal2 s 112782 -960 112894 480 0 FreeSans 448 90 0 0 wbs_dat_i[28]
port 595 nsew signal input
flabel metal2 s 116370 -960 116482 480 0 FreeSans 448 90 0 0 wbs_dat_i[29]
port 596 nsew signal input
flabel metal2 s 18206 -960 18318 480 0 FreeSans 448 90 0 0 wbs_dat_i[2]
port 597 nsew signal input
flabel metal2 s 119866 -960 119978 480 0 FreeSans 448 90 0 0 wbs_dat_i[30]
port 598 nsew signal input
flabel metal2 s 123454 -960 123566 480 0 FreeSans 448 90 0 0 wbs_dat_i[31]
port 599 nsew signal input
flabel metal2 s 22990 -960 23102 480 0 FreeSans 448 90 0 0 wbs_dat_i[3]
port 600 nsew signal input
flabel metal2 s 27682 -960 27794 480 0 FreeSans 448 90 0 0 wbs_dat_i[4]
port 601 nsew signal input
flabel metal2 s 31270 -960 31382 480 0 FreeSans 448 90 0 0 wbs_dat_i[5]
port 602 nsew signal input
flabel metal2 s 34766 -960 34878 480 0 FreeSans 448 90 0 0 wbs_dat_i[6]
port 603 nsew signal input
flabel metal2 s 38354 -960 38466 480 0 FreeSans 448 90 0 0 wbs_dat_i[7]
port 604 nsew signal input
flabel metal2 s 41850 -960 41962 480 0 FreeSans 448 90 0 0 wbs_dat_i[8]
port 605 nsew signal input
flabel metal2 s 45438 -960 45550 480 0 FreeSans 448 90 0 0 wbs_dat_i[9]
port 606 nsew signal input
flabel metal2 s 9926 -960 10038 480 0 FreeSans 448 90 0 0 wbs_dat_o[0]
port 607 nsew signal tristate
flabel metal2 s 50130 -960 50242 480 0 FreeSans 448 90 0 0 wbs_dat_o[10]
port 608 nsew signal tristate
flabel metal2 s 53718 -960 53830 480 0 FreeSans 448 90 0 0 wbs_dat_o[11]
port 609 nsew signal tristate
flabel metal2 s 57214 -960 57326 480 0 FreeSans 448 90 0 0 wbs_dat_o[12]
port 610 nsew signal tristate
flabel metal2 s 60802 -960 60914 480 0 FreeSans 448 90 0 0 wbs_dat_o[13]
port 611 nsew signal tristate
flabel metal2 s 64298 -960 64410 480 0 FreeSans 448 90 0 0 wbs_dat_o[14]
port 612 nsew signal tristate
flabel metal2 s 67886 -960 67998 480 0 FreeSans 448 90 0 0 wbs_dat_o[15]
port 613 nsew signal tristate
flabel metal2 s 71474 -960 71586 480 0 FreeSans 448 90 0 0 wbs_dat_o[16]
port 614 nsew signal tristate
flabel metal2 s 74970 -960 75082 480 0 FreeSans 448 90 0 0 wbs_dat_o[17]
port 615 nsew signal tristate
flabel metal2 s 78558 -960 78670 480 0 FreeSans 448 90 0 0 wbs_dat_o[18]
port 616 nsew signal tristate
flabel metal2 s 82054 -960 82166 480 0 FreeSans 448 90 0 0 wbs_dat_o[19]
port 617 nsew signal tristate
flabel metal2 s 14710 -960 14822 480 0 FreeSans 448 90 0 0 wbs_dat_o[1]
port 618 nsew signal tristate
flabel metal2 s 85642 -960 85754 480 0 FreeSans 448 90 0 0 wbs_dat_o[20]
port 619 nsew signal tristate
flabel metal2 s 89138 -960 89250 480 0 FreeSans 448 90 0 0 wbs_dat_o[21]
port 620 nsew signal tristate
flabel metal2 s 92726 -960 92838 480 0 FreeSans 448 90 0 0 wbs_dat_o[22]
port 621 nsew signal tristate
flabel metal2 s 96222 -960 96334 480 0 FreeSans 448 90 0 0 wbs_dat_o[23]
port 622 nsew signal tristate
flabel metal2 s 99810 -960 99922 480 0 FreeSans 448 90 0 0 wbs_dat_o[24]
port 623 nsew signal tristate
flabel metal2 s 103306 -960 103418 480 0 FreeSans 448 90 0 0 wbs_dat_o[25]
port 624 nsew signal tristate
flabel metal2 s 106894 -960 107006 480 0 FreeSans 448 90 0 0 wbs_dat_o[26]
port 625 nsew signal tristate
flabel metal2 s 110482 -960 110594 480 0 FreeSans 448 90 0 0 wbs_dat_o[27]
port 626 nsew signal tristate
flabel metal2 s 113978 -960 114090 480 0 FreeSans 448 90 0 0 wbs_dat_o[28]
port 627 nsew signal tristate
flabel metal2 s 117566 -960 117678 480 0 FreeSans 448 90 0 0 wbs_dat_o[29]
port 628 nsew signal tristate
flabel metal2 s 19402 -960 19514 480 0 FreeSans 448 90 0 0 wbs_dat_o[2]
port 629 nsew signal tristate
flabel metal2 s 121062 -960 121174 480 0 FreeSans 448 90 0 0 wbs_dat_o[30]
port 630 nsew signal tristate
flabel metal2 s 124650 -960 124762 480 0 FreeSans 448 90 0 0 wbs_dat_o[31]
port 631 nsew signal tristate
flabel metal2 s 24186 -960 24298 480 0 FreeSans 448 90 0 0 wbs_dat_o[3]
port 632 nsew signal tristate
flabel metal2 s 28878 -960 28990 480 0 FreeSans 448 90 0 0 wbs_dat_o[4]
port 633 nsew signal tristate
flabel metal2 s 32374 -960 32486 480 0 FreeSans 448 90 0 0 wbs_dat_o[5]
port 634 nsew signal tristate
flabel metal2 s 35962 -960 36074 480 0 FreeSans 448 90 0 0 wbs_dat_o[6]
port 635 nsew signal tristate
flabel metal2 s 39550 -960 39662 480 0 FreeSans 448 90 0 0 wbs_dat_o[7]
port 636 nsew signal tristate
flabel metal2 s 43046 -960 43158 480 0 FreeSans 448 90 0 0 wbs_dat_o[8]
port 637 nsew signal tristate
flabel metal2 s 46634 -960 46746 480 0 FreeSans 448 90 0 0 wbs_dat_o[9]
port 638 nsew signal tristate
flabel metal2 s 11122 -960 11234 480 0 FreeSans 448 90 0 0 wbs_sel_i[0]
port 639 nsew signal input
flabel metal2 s 15906 -960 16018 480 0 FreeSans 448 90 0 0 wbs_sel_i[1]
port 640 nsew signal input
flabel metal2 s 20598 -960 20710 480 0 FreeSans 448 90 0 0 wbs_sel_i[2]
port 641 nsew signal input
flabel metal2 s 25290 -960 25402 480 0 FreeSans 448 90 0 0 wbs_sel_i[3]
port 642 nsew signal input
flabel metal2 s 5234 -960 5346 480 0 FreeSans 448 90 0 0 wbs_stb_i
port 643 nsew signal input
flabel metal2 s 6430 -960 6542 480 0 FreeSans 448 90 0 0 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
